* NGSPICE file created from heichips25_tiny_wrapper2.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_1 abstract view
.subckt sg13g2_dfrbpq_1 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_nand4_1 abstract view
.subckt sg13g2_nand4_1 B C A Y VDD VSS D
.ends

* Black-box entry subcircuit for sg13g2_tielo abstract view
.subckt sg13g2_tielo VDD VSS L_LO
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xor2_1 abstract view
.subckt sg13g2_xor2_1 B A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_1 abstract view
.subckt sg13g2_nor2b_1 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tiehi abstract view
.subckt sg13g2_tiehi VDD VSS L_HI
.ends

* Black-box entry subcircuit for sg13g2_dlygate4sd3_1 abstract view
.subckt sg13g2_dlygate4sd3_1 A VDD VSS X
.ends

* Black-box entry subcircuit for sg13g2_a22oi_1 abstract view
.subckt sg13g2_a22oi_1 Y B1 B2 A2 A1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor3_1 abstract view
.subckt sg13g2_nor3_1 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux2_1 abstract view
.subckt sg13g2_mux2_1 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xnor2_1 abstract view
.subckt sg13g2_xnor2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_16 abstract view
.subckt sg13g2_buf_16 X A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a221oi_1 abstract view
.subckt sg13g2_a221oi_1 VDD VSS B2 C1 B1 A1 Y A2
.ends

* Black-box entry subcircuit for sg13g2_and2_1 abstract view
.subckt sg13g2_and2_1 A B X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and3_1 abstract view
.subckt sg13g2_and3_1 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3b_1 abstract view
.subckt sg13g2_nand3b_1 B C Y VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_nand3_1 abstract view
.subckt sg13g2_nand3_1 B C A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21o_1 abstract view
.subckt sg13g2_a21o_1 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor4_1 abstract view
.subckt sg13g2_nor4_1 A B C D Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and4_1 abstract view
.subckt sg13g2_and4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or4_1 abstract view
.subckt sg13g2_or4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_2 abstract view
.subckt sg13g2_buf_2 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux4_1 abstract view
.subckt sg13g2_mux4_1 S0 A0 A1 A2 A3 S1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or3_1 abstract view
.subckt sg13g2_or3_1 A B C X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_4 abstract view
.subckt sg13g2_inv_4 A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor4_2 abstract view
.subckt sg13g2_nor4_2 A B C Y VSS VDD D
.ends

* Black-box entry subcircuit for sg13g2_inv_2 abstract view
.subckt sg13g2_inv_2 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_4 abstract view
.subckt sg13g2_buf_4 X A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_lgcp_1 abstract view
.subckt sg13g2_lgcp_1 GATE CLK GCLK VDD VSS
.ends

.subckt heichips25_tiny_wrapper2 VGND VPWR clk ena rst_n ui_in[0] ui_in[1] ui_in[2]
+ ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3]
+ uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3]
+ uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3]
+ uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3]
+ uo_out[4] uo_out[5] uo_out[6] uo_out[7]
XFILLER_36_19 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2823_ net560 VGND VPWR heichips25_can_lehmann_fsm/_0048_
+ heichips25_can_lehmann_fsm__2823_/Q clknet_leaf_9_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2754_ heichips25_can_lehmann_fsm/net498 VPWR heichips25_can_lehmann_fsm/_0843_
+ VGND heichips25_can_lehmann_fsm__3052_/Q heichips25_can_lehmann_fsm/net426 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__1705_ heichips25_can_lehmann_fsm/_1029_ heichips25_can_lehmann_fsm/_1028_
+ heichips25_can_lehmann_fsm/_1022_ VPWR VGND sg13g2_nand2b_1
XFILLER_23_612 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2685_ VGND VPWR heichips25_can_lehmann_fsm/_0874_ heichips25_can_lehmann_fsm/net359
+ heichips25_can_lehmann_fsm/_0242_ heichips25_can_lehmann_fsm/_0808_ sg13g2_a21oi_1
Xclkbuf_4_12_0_heichips25_sap3\_sap_3_inst.alu_inst.clk clknet_0_heichips25_sap3\/sap_3_inst.alu_inst.clk
+ clknet_4_12_0_heichips25_sap3\/sap_3_inst.alu_inst.clk VPWR VGND sg13g2_buf_8
Xheichips25_can_lehmann_fsm__1636_ VPWR heichips25_can_lehmann_fsm/_0960_ heichips25_can_lehmann_fsm/net965
+ VGND sg13g2_inv_1
XFILLER_23_667 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1567_ VPWR heichips25_can_lehmann_fsm/_0891_ heichips25_can_lehmann_fsm/net889
+ VGND sg13g2_inv_1
XFILLER_7_7 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2119_ heichips25_can_lehmann_fsm/_0455_ heichips25_can_lehmann_fsm/_0456_
+ heichips25_can_lehmann_fsm/_0454_ heichips25_can_lehmann_fsm/_0458_ VPWR VGND heichips25_can_lehmann_fsm/_0457_
+ sg13g2_nand4_1
XFILLER_45_214 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3120_ heichips25_sap3/_1581_ VPWR heichips25_sap3/_0733_ VGND heichips25_sap3/net243
+ heichips25_sap3/_0307_ sg13g2_o21ai_1
XFILLER_26_41 VPWR VGND sg13g2_fill_2
X_16__518 VPWR VGND net517 sg13g2_tielo
Xheichips25_sap3__3051_ heichips25_sap3/_0664_ heichips25_sap3/_0660_ heichips25_sap3/_0662_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__2002_ VPWR heichips25_sap3/_1428_ heichips25_sap3__4040_/Q VGND
+ sg13g2_inv_1
XFILLER_42_51 VPWR VGND sg13g2_fill_2
XFILLER_9_126 VPWR VGND sg13g2_decap_8
XFILLER_9_137 VPWR VGND sg13g2_decap_4
XFILLER_10_840 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3953_ heichips25_sap3/net440 VGND VPWR heichips25_sap3/_0094_ heichips25_sap3__3953_/Q
+ heichips25_sap3__4017_/CLK sg13g2_dfrbpq_1
Xheichips25_sap3__3884_ heichips25_sap3/net450 VGND VPWR heichips25_sap3/_0025_ heichips25_sap3__3884_/Q
+ heichips25_sap3__3922_/CLK sg13g2_dfrbpq_1
Xheichips25_sap3__2904_ heichips25_sap3/_0540_ heichips25_sap3/_0541_ heichips25_sap3/_0539_
+ heichips25_sap3/_0544_ VPWR VGND heichips25_sap3/_0543_ sg13g2_nand4_1
Xheichips25_sap3__2835_ heichips25_sap3/net159 VPWR heichips25_sap3/_0478_ VGND heichips25_sap3/net284
+ heichips25_sap3__3917_/Q sg13g2_o21ai_1
Xheichips25_sap3__2766_ heichips25_sap3/_0411_ heichips25_sap3/_0381_ heichips25_sap3/_0412_
+ VPWR VGND sg13g2_xor2_1
XFILLER_1_571 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2697_ heichips25_sap3/_1887_ heichips25_sap3/_1894_ heichips25_sap3/_0343_
+ VPWR VGND sg13g2_nor2b_1
Xheichips25_sap3__3318_ heichips25_sap3/_0929_ heichips25_sap3/net97 heichips25_sap3/_0928_
+ VPWR VGND sg13g2_nand2_1
XFILLER_45_792 VPWR VGND sg13g2_fill_2
XFILLER_17_461 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3249_ heichips25_sap3/_0731_ heichips25_sap3/net166 heichips25_sap3/_0862_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_can_lehmann_fsm__2470_ heichips25_can_lehmann_fsm/net487 VPWR heichips25_can_lehmann_fsm/_0701_
+ VGND heichips25_can_lehmann_fsm__2910_/Q heichips25_can_lehmann_fsm/net418 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__3022_ net706 VGND VPWR heichips25_can_lehmann_fsm/_0247_
+ heichips25_can_lehmann_fsm__3022_/Q clknet_leaf_6_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2870__756 VPWR VGND net755 sg13g2_tiehi
XFILLER_28_748 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2806_ net594 VGND VPWR heichips25_can_lehmann_fsm/net1237
+ heichips25_can_lehmann_fsm__2806_/Q clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_42_217 VPWR VGND sg13g2_decap_8
XFILLER_27_269 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2737_ VGND VPWR heichips25_can_lehmann_fsm/_0861_ heichips25_can_lehmann_fsm/net390
+ heichips25_can_lehmann_fsm/_0268_ heichips25_can_lehmann_fsm/_0834_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2668_ heichips25_can_lehmann_fsm/net483 VPWR heichips25_can_lehmann_fsm/_0800_
+ VGND heichips25_can_lehmann_fsm__3008_/Q heichips25_can_lehmann_fsm/net375 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm_hold858 heichips25_can_lehmann_fsm__2850_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net857 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__1619_ VPWR heichips25_can_lehmann_fsm/_0943_ heichips25_can_lehmann_fsm/net916
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm_hold847 heichips25_can_lehmann_fsm__2975_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net846 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold869 heichips25_can_lehmann_fsm/_0234_ VPWR VGND heichips25_can_lehmann_fsm/net868
+ sg13g2_dlygate4sd3_1
XFILLER_12_21 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2599_ VGND VPWR heichips25_can_lehmann_fsm/_0898_ heichips25_can_lehmann_fsm/net407
+ heichips25_can_lehmann_fsm/_0199_ heichips25_can_lehmann_fsm/_0765_ sg13g2_a21oi_1
XFILLER_10_169 VPWR VGND sg13g2_decap_4
XFILLER_12_76 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2620_ heichips25_sap3/_0289_ heichips25_sap3/net1130 heichips25_sap3/_1431_
+ VPWR VGND sg13g2_nand2_1
XFILLER_5_4 VPWR VGND sg13g2_decap_8
XFILLER_2_324 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2916__664 VPWR VGND net663 sg13g2_tiehi
Xheichips25_sap3__2551_ heichips25_sap3/_0226_ heichips25_sap3/net80 heichips25_sap3__4022_/Q
+ heichips25_sap3/net85 heichips25_sap3__3950_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2482_ heichips25_sap3/_1883_ heichips25_sap3/_1884_ heichips25_sap3/net168
+ heichips25_sap3/_1895_ VPWR VGND sg13g2_nor3_1
XFILLER_18_225 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3103_ heichips25_sap3/_0716_ heichips25_sap3/_0654_ heichips25_sap3/_1441_
+ heichips25_sap3/_1467_ heichips25_sap3/_1457_ VPWR VGND sg13g2_a22oi_1
XFILLER_14_431 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3034_ heichips25_sap3/net263 VPWR heichips25_sap3/_0647_ VGND heichips25_sap3/_0644_
+ heichips25_sap3/_0645_ sg13g2_o21ai_1
XFILLER_14_464 VPWR VGND sg13g2_fill_2
XFILLER_18_1015 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3936_ heichips25_sap3/net441 VGND VPWR heichips25_sap3/_0077_ heichips25_sap3__3936_/Q
+ heichips25_sap3__4016_/CLK sg13g2_dfrbpq_1
XFILLER_6_674 VPWR VGND sg13g2_fill_2
XFILLER_5_162 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3867_ heichips25_sap3__3886_/Q heichips25_sap3/net1143 heichips25_sap3/_0007_
+ heichips25_sap3/_0194_ VPWR VGND sg13g2_mux2_1
Xheichips25_sap3__2818_ heichips25_sap3/_0462_ heichips25_sap3/_1381_ heichips25_sap3/net212
+ VPWR VGND sg13g2_xnor2_1
Xheichips25_sap3__3798_ heichips25_sap3/_1307_ heichips25_sap3/_1278_ heichips25_sap3__4006_/Q
+ heichips25_sap3/_1265_ heichips25_sap3__3998_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2817__573 VPWR VGND net572 sg13g2_tiehi
Xheichips25_sap3__2749_ heichips25_sap3/_1383_ heichips25_sap3__3919_/Q heichips25_sap3/_0395_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_can_lehmann_fsm__1970_ VGND VPWR heichips25_can_lehmann_fsm/_0330_ heichips25_can_lehmann_fsm/_0329_
+ heichips25_can_lehmann_fsm/net192 sg13g2_or2_1
XFILLER_49_361 VPWR VGND sg13g2_decap_8
XFILLER_37_578 VPWR VGND sg13g2_fill_2
XFILLER_18_792 VPWR VGND sg13g2_decap_8
XFILLER_24_228 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2522_ heichips25_can_lehmann_fsm/net483 VPWR heichips25_can_lehmann_fsm/_0727_
+ VGND heichips25_can_lehmann_fsm/net1079 heichips25_can_lehmann_fsm/net415 sg13g2_o21ai_1
XFILLER_33_751 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2453_ VGND VPWR heichips25_can_lehmann_fsm/_0934_ heichips25_can_lehmann_fsm/net365
+ heichips25_can_lehmann_fsm/_0126_ heichips25_can_lehmann_fsm/_0692_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2384_ heichips25_can_lehmann_fsm/net481 VPWR heichips25_can_lehmann_fsm/_0658_
+ VGND heichips25_can_lehmann_fsm/net912 heichips25_can_lehmann_fsm/net372 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm_fanout500 heichips25_can_lehmann_fsm/net502 heichips25_can_lehmann_fsm/net500
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm__3005_ net553 VGND VPWR heichips25_can_lehmann_fsm/_0230_
+ heichips25_can_lehmann_fsm__3005_/Q clknet_leaf_12_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__3046__663 VPWR VGND net662 sg13g2_tiehi
XFILLER_43_559 VPWR VGND sg13g2_decap_8
XFILLER_15_228 VPWR VGND sg13g2_fill_1
XFILLER_15_239 VPWR VGND sg13g2_fill_2
XFILLER_7_416 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__1982_ VPWR heichips25_sap3/_1408_ heichips25_sap3__3984_/Q VGND
+ sg13g2_inv_1
Xheichips25_sap3__3721_ heichips25_sap3__4022_/Q heichips25_sap3/_1068_ heichips25_sap3/net117
+ heichips25_sap3/_0163_ VPWR VGND sg13g2_mux2_1
Xheichips25_can_lehmann_fsm__2957__797 VPWR VGND net796 sg13g2_tiehi
Xheichips25_sap3__3652_ heichips25_sap3/_1199_ VPWR heichips25_sap3/_1200_ VGND heichips25_sap3/net48
+ heichips25_sap3/net51 sg13g2_o21ai_1
Xheichips25_sap3__2603_ heichips25_sap3/_0275_ heichips25_sap3/_0273_ heichips25_sap3/_0274_
+ VPWR VGND sg13g2_xnor2_1
Xheichips25_sap3__3583_ heichips25_sap3__3967_/Q heichips25_sap3/net135 heichips25_sap3/_1160_
+ VPWR VGND sg13g2_nor2_1
XFILLER_38_309 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2534_ VGND VPWR heichips25_sap3/_0206_ heichips25_sap3/_0210_ heichips25_sap3/_0211_
+ heichips25_sap3/net67 sg13g2_a21oi_1
XFILLER_19_501 VPWR VGND sg13g2_fill_2
XFILLER_19_512 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2465_ heichips25_sap3/net215 heichips25_sap3/_1877_ heichips25_sap3/_1878_
+ VPWR VGND sg13g2_nor2_1
Xclkbuf_5_19__f_heichips25_sap3\_sap_3_inst.alu_inst.clk clkload24/A clknet_4_9_0_heichips25_sap3\/sap_3_inst.alu_inst.clk
+ VPWR VGND sg13g2_buf_16
Xheichips25_sap3__2396_ heichips25_sap3/_1815_ heichips25_sap3/net155 heichips25_sap3/_1814_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__4066_ heichips25_sap3/net433 VGND VPWR heichips25_sap3/_0006_ heichips25_sap3__4066_/Q
+ net825 sg13g2_dfrbpq_1
Xheichips25_sap3__3017_ heichips25_sap3/_0634_ VPWR heichips25_sap3/_0067_ VGND heichips25_sap3/net232
+ heichips25_sap3/_0242_ sg13g2_o21ai_1
XFILLER_15_784 VPWR VGND sg13g2_fill_1
XFILLER_14_294 VPWR VGND sg13g2_decap_4
XFILLER_9_99 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3919_ heichips25_sap3/net448 VGND VPWR heichips25_sap3/_0060_ heichips25_sap3__3919_/Q
+ heichips25_sap3__3920_/CLK sg13g2_dfrbpq_1
XFILLER_29_309 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__1953_ VPWR VGND heichips25_can_lehmann_fsm/net195 heichips25_can_lehmann_fsm/_0315_
+ heichips25_can_lehmann_fsm/_0314_ heichips25_can_lehmann_fsm/_0308_ heichips25_can_lehmann_fsm/_0003_
+ heichips25_can_lehmann_fsm/_0311_ sg13g2_a221oi_1
XFILLER_38_898 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1884_ heichips25_can_lehmann_fsm/_1197_ heichips25_can_lehmann_fsm/net338
+ heichips25_can_lehmann_fsm/_1165_ heichips25_can_lehmann_fsm/_1198_ VPWR VGND sg13g2_mux2_1
Xheichips25_sap3_fanout437 _01_ heichips25_sap3/net437 VPWR VGND sg13g2_buf_1
Xheichips25_sap3_fanout448 heichips25_sap3/net449 heichips25_sap3/net448 VPWR VGND
+ sg13g2_buf_1
XFILLER_25_559 VPWR VGND sg13g2_decap_8
Xheichips25_sap3_fanout459 heichips25_sap3/net461 heichips25_sap3/net459 VPWR VGND
+ sg13g2_buf_1
XFILLER_40_507 VPWR VGND sg13g2_fill_2
Xheichips25_sap3_hold1059 heichips25_sap3__4073_/A VPWR VGND heichips25_sap3/net1058
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__2505_ VGND VPWR heichips25_can_lehmann_fsm/_0921_ heichips25_can_lehmann_fsm/net366
+ heichips25_can_lehmann_fsm/_0152_ heichips25_can_lehmann_fsm/_0718_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2436_ heichips25_can_lehmann_fsm/net477 VPWR heichips25_can_lehmann_fsm/_0684_
+ VGND heichips25_can_lehmann_fsm/net989 heichips25_can_lehmann_fsm/net368 sg13g2_o21ai_1
XFILLER_20_264 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2367_ VGND VPWR heichips25_can_lehmann_fsm/_0960_ heichips25_can_lehmann_fsm/net431
+ heichips25_can_lehmann_fsm/_0083_ heichips25_can_lehmann_fsm/_0649_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2298_ heichips25_can_lehmann_fsm/_0609_ heichips25_can_lehmann_fsm/net1200
+ heichips25_can_lehmann_fsm/_0608_ VPWR VGND sg13g2_xnor2_1
Xheichips25_can_lehmann_fsm_fanout330 heichips25_can_lehmann_fsm/_1175_ heichips25_can_lehmann_fsm/net330
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout363 heichips25_can_lehmann_fsm/net364 heichips25_can_lehmann_fsm/net363
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout374 heichips25_can_lehmann_fsm/net375 heichips25_can_lehmann_fsm/net374
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout352 heichips25_can_lehmann_fsm/net1273 heichips25_can_lehmann_fsm/net352
+ VPWR VGND sg13g2_buf_1
XFILLER_0_625 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_fanout396 heichips25_can_lehmann_fsm/net397 heichips25_can_lehmann_fsm/net396
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout385 heichips25_can_lehmann_fsm/net387 heichips25_can_lehmann_fsm/net385
+ VPWR VGND sg13g2_buf_1
Xheichips25_sap3__2250_ heichips25_sap3/_1462_ heichips25_sap3/_1615_ heichips25_sap3/_1655_
+ heichips25_sap3/_1671_ VPWR VGND sg13g2_nor3_1
XFILLER_16_504 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2181_ heichips25_sap3/_1602_ heichips25_sap3/_1551_ heichips25_sap3/_1567_
+ VPWR VGND sg13g2_nand2_1
XFILLER_16_526 VPWR VGND sg13g2_fill_2
XFILLER_18_97 VPWR VGND sg13g2_fill_2
XFILLER_43_367 VPWR VGND sg13g2_fill_2
XFILLER_12_754 VPWR VGND sg13g2_decap_4
XFILLER_7_257 VPWR VGND sg13g2_decap_4
XFILLER_3_430 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__1965_ VPWR heichips25_sap3/_1391_ heichips25_sap3__3948_/Q VGND
+ sg13g2_inv_1
XFILLER_4_964 VPWR VGND sg13g2_fill_2
XFILLER_3_463 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3704_ VGND VPWR heichips25_sap3/_1100_ heichips25_sap3/_1204_ heichips25_sap3/_1235_
+ heichips25_sap3/net115 sg13g2_a21oi_1
XFILLER_3_485 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3635_ heichips25_sap3/_1190_ VPWR heichips25_sap3/_0129_ VGND heichips25_sap3/_1063_
+ heichips25_sap3/net93 sg13g2_o21ai_1
Xheichips25_sap3__3566_ heichips25_sap3/net134 heichips25_sap3/_1054_ heichips25_sap3/_1147_
+ VPWR VGND sg13g2_nor2_1
XFILLER_15_6 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3497_ heichips25_sap3/net97 heichips25_sap3/_0911_ heichips25_sap3/_1093_
+ VPWR VGND sg13g2_and2_1
Xheichips25_sap3__2517_ heichips25_sap3/_1928_ heichips25_sap3/net82 heichips25_sap3__3963_/Q
+ heichips25_sap3/net88 heichips25_sap3__3939_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2448_ heichips25_sap3/_1863_ heichips25_sap3/_1860_ heichips25_sap3/_1861_
+ heichips25_sap3/_1862_ VPWR VGND sg13g2_and3_1
Xheichips25_sap3__2379_ VGND VPWR heichips25_sap3/_1795_ heichips25_sap3/_1799_ heichips25_sap3/_1800_
+ heichips25_sap3/net66 sg13g2_a21oi_1
Xheichips25_sap3__4049_ heichips25_sap3/net451 VGND VPWR heichips25_sap3/_0190_ heichips25_sap3__4049_/Q
+ clknet_leaf_23_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2221_ heichips25_can_lehmann_fsm/net1217 VPWR heichips25_can_lehmann_fsm/_0547_
+ VGND heichips25_can_lehmann_fsm/net1279 heichips25_can_lehmann_fsm/_1104_ sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2152_ VGND VPWR heichips25_can_lehmann_fsm/_1162_ heichips25_can_lehmann_fsm/_0482_
+ heichips25_can_lehmann_fsm/_0491_ heichips25_can_lehmann_fsm/_1139_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2083_ VPWR VGND heichips25_can_lehmann_fsm__2799_/Q heichips25_can_lehmann_fsm/net182
+ heichips25_can_lehmann_fsm/net190 net15 heichips25_can_lehmann_fsm/_0426_ heichips25_can_lehmann_fsm/net195
+ sg13g2_a221oi_1
XFILLER_29_106 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2985_ net684 VGND VPWR heichips25_can_lehmann_fsm/_0210_
+ heichips25_can_lehmann_fsm__2985_/Q clknet_leaf_16_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1936_ heichips25_can_lehmann_fsm/_0296_ heichips25_can_lehmann_fsm/_0297_
+ heichips25_can_lehmann_fsm/_0295_ heichips25_can_lehmann_fsm/_0299_ VPWR VGND heichips25_can_lehmann_fsm/_0298_
+ sg13g2_nand4_1
Xheichips25_sap3_fanout212 heichips25_sap3/_1889_ heichips25_sap3/net212 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout201 heichips25_sap3/_0624_ heichips25_sap3/net201 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout223 heichips25_sap3/_1622_ heichips25_sap3/net223 VPWR VGND
+ sg13g2_buf_1
Xheichips25_can_lehmann_fsm__1867_ heichips25_can_lehmann_fsm/_1179_ heichips25_can_lehmann_fsm/_1180_
+ heichips25_can_lehmann_fsm/_1178_ heichips25_can_lehmann_fsm/_1182_ VPWR VGND heichips25_can_lehmann_fsm/_1181_
+ sg13g2_nand4_1
Xheichips25_sap3_fanout256 heichips25_sap3/_1442_ heichips25_sap3/net256 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout245 heichips25_sap3/_1509_ heichips25_sap3/net245 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout234 heichips25_sap3/net235 heichips25_sap3/net234 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout267 heichips25_sap3__3925_/Q heichips25_sap3/net267 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout278 heichips25_sap3/net279 heichips25_sap3/net278 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout289 heichips25_sap3__3899_/Q heichips25_sap3/net289 VPWR VGND
+ sg13g2_buf_1
Xheichips25_can_lehmann_fsm__1798_ heichips25_can_lehmann_fsm/_1114_ heichips25_can_lehmann_fsm/_1111_
+ heichips25_can_lehmann_fsm/_1113_ heichips25_can_lehmann_fsm/net301 heichips25_can_lehmann_fsm/_0949_
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2419_ VGND VPWR heichips25_can_lehmann_fsm/_0944_ heichips25_can_lehmann_fsm/net384
+ heichips25_can_lehmann_fsm/_0109_ heichips25_can_lehmann_fsm/_0675_ sg13g2_a21oi_1
XFILLER_5_728 VPWR VGND sg13g2_fill_2
XFILLER_4_227 VPWR VGND sg13g2_decap_8
XFILLER_20_21 VPWR VGND sg13g2_decap_8
XFILLER_1_912 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm_fanout182 heichips25_can_lehmann_fsm/net183 heichips25_can_lehmann_fsm/net182
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout160 heichips25_can_lehmann_fsm/net163 heichips25_can_lehmann_fsm/net160
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout171 heichips25_can_lehmann_fsm/net173 heichips25_can_lehmann_fsm/net171
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout193 heichips25_can_lehmann_fsm/net194 heichips25_can_lehmann_fsm/net193
+ VPWR VGND sg13g2_buf_1
Xheichips25_sap3__3420_ VGND VPWR heichips25_sap3/net126 heichips25_sap3/_1024_ heichips25_sap3/_1027_
+ heichips25_sap3/_1026_ sg13g2_a21oi_1
XFILLER_1_989 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3351_ heichips25_sap3/_0960_ heichips25_sap3__3959_/Q heichips25_sap3/net144
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__2302_ heichips25_sap3/net234 heichips25_sap3/_1722_ heichips25_sap3/_1723_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__3282_ heichips25_sap3/_0894_ heichips25_sap3/net123 heichips25_sap3/_0893_
+ VPWR VGND sg13g2_nand2_1
XFILLER_28_150 VPWR VGND sg13g2_decap_8
XFILLER_45_40 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2233_ heichips25_sap3/_1653_ heichips25_sap3/net67 heichips25_sap3/_1654_
+ VPWR VGND heichips25_sap3/_1650_ sg13g2_nand3b_1
XFILLER_17_835 VPWR VGND sg13g2_fill_1
XFILLER_45_73 VPWR VGND sg13g2_decap_8
XFILLER_16_345 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2164_ heichips25_sap3/_1585_ heichips25_sap3/_1576_ heichips25_sap3/net243
+ heichips25_sap3/_1563_ heichips25_sap3/net242 VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2095_ heichips25_sap3/_1445_ heichips25_sap3/_1505_ heichips25_sap3/_1365_
+ heichips25_sap3/_1516_ VPWR VGND sg13g2_nand3_1
XFILLER_31_359 VPWR VGND sg13g2_fill_1
XFILLER_40_882 VPWR VGND sg13g2_fill_2
XFILLER_8_555 VPWR VGND sg13g2_fill_2
XFILLER_6_34 VPWR VGND sg13g2_decap_8
XFILLER_8_588 VPWR VGND sg13g2_decap_8
XFILLER_6_67 VPWR VGND sg13g2_fill_1
XFILLER_6_89 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2997_ VGND VPWR heichips25_sap3/_0212_ heichips25_sap3/net201 heichips25_sap3/_0056_
+ heichips25_sap3/_0625_ sg13g2_a21oi_1
Xheichips25_sap3__1948_ VPWR heichips25_sap3/_1374_ heichips25_sap3/net274 VGND sg13g2_inv_1
XFILLER_20_4 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3618_ heichips25_sap3/net141 heichips25_sap3/_1064_ heichips25_sap3/_1181_
+ VPWR VGND sg13g2_and2_1
Xheichips25_sap3__3549_ heichips25_sap3/_1136_ VPWR heichips25_sap3/_0097_ VGND heichips25_sap3/_1390_
+ heichips25_sap3/net56 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2770_ heichips25_can_lehmann_fsm/net481 VPWR heichips25_can_lehmann_fsm/_0851_
+ VGND heichips25_can_lehmann_fsm/net1137 heichips25_can_lehmann_fsm/net400 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__1721_ uo_out_fsm\[2\] heichips25_can_lehmann_fsm/_1041_
+ heichips25_can_lehmann_fsm/_1042_ VPWR VGND sg13g2_nand2_1
Xheichips25_can_lehmann_fsm__1652_ VPWR heichips25_can_lehmann_fsm/_0976_ heichips25_can_lehmann_fsm__2797_/Q
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__1583_ VPWR heichips25_can_lehmann_fsm/_0907_ heichips25_can_lehmann_fsm/net1027
+ VGND sg13g2_inv_1
Xclkbuf_5_2__f_heichips25_sap3\_sap_3_inst.alu_inst.clk heichips25_sap3__4014_/CLK
+ clknet_4_1_0_heichips25_sap3\/sap_3_inst.alu_inst.clk VPWR VGND sg13g2_buf_16
Xheichips25_can_lehmann_fsm__2204_ heichips25_can_lehmann_fsm/_0534_ heichips25_can_lehmann_fsm/net1180
+ heichips25_can_lehmann_fsm/_1102_ VPWR VGND sg13g2_xnor2_1
Xheichips25_can_lehmann_fsm__2135_ VGND VPWR heichips25_can_lehmann_fsm/_0942_ heichips25_can_lehmann_fsm/net303
+ heichips25_can_lehmann_fsm/_0474_ heichips25_can_lehmann_fsm/_0473_ sg13g2_a21oi_1
XFILLER_44_1000 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2066_ VPWR VGND heichips25_can_lehmann_fsm/_0977_ heichips25_can_lehmann_fsm/net181
+ heichips25_can_lehmann_fsm/net184 heichips25_can_lehmann_fsm/net347 heichips25_can_lehmann_fsm/_0413_
+ heichips25_can_lehmann_fsm/net188 sg13g2_a221oi_1
XFILLER_39_971 VPWR VGND sg13g2_fill_1
XFILLER_38_492 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2968_ net752 VGND VPWR heichips25_can_lehmann_fsm/_0193_
+ heichips25_can_lehmann_fsm__2968_/Q clknet_leaf_20_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2899_ net697 VGND VPWR heichips25_can_lehmann_fsm/net1057
+ heichips25_can_lehmann_fsm__2899_/Q clknet_leaf_21_clk sg13g2_dfrbpq_1
XFILLER_25_131 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1919_ VPWR heichips25_can_lehmann_fsm/_1232_ heichips25_can_lehmann_fsm/_1231_
+ VGND sg13g2_inv_1
XFILLER_14_838 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2880__736 VPWR VGND net735 sg13g2_tiehi
Xheichips25_can_lehmann_fsm_hold1110 heichips25_can_lehmann_fsm__2958_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1109 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1154 heichips25_can_lehmann_fsm__3027_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1153 sg13g2_dlygate4sd3_1
XFILLER_9_308 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm_hold1165 heichips25_can_lehmann_fsm__3036_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1164 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1143 heichips25_can_lehmann_fsm__3057_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1142 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1187 heichips25_can_lehmann_fsm__2813_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1186 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1176 heichips25_can_lehmann_fsm/_0044_ VPWR VGND heichips25_can_lehmann_fsm/net1175
+ sg13g2_dlygate4sd3_1
Xheichips25_sap3__2920_ heichips25_sap3/net69 heichips25_sap3/net279 heichips25_sap3/_0559_
+ heichips25_sap3/_0045_ VPWR VGND sg13g2_a21o_1
XFILLER_31_53 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2851_ VGND VPWR heichips25_sap3/_0375_ heichips25_sap3/net64 heichips25_sap3/_0494_
+ heichips25_sap3/net204 sg13g2_a21oi_1
XFILLER_31_64 VPWR VGND sg13g2_fill_2
XFILLER_5_558 VPWR VGND sg13g2_fill_2
Xheichips25_sap3_fanout62 heichips25_sap3/_0829_ heichips25_sap3/net62 VPWR VGND sg13g2_buf_1
Xheichips25_sap3_fanout51 heichips25_sap3/_0898_ heichips25_sap3/net51 VPWR VGND sg13g2_buf_1
Xheichips25_sap3_fanout84 heichips25_sap3/_1739_ heichips25_sap3/net84 VPWR VGND sg13g2_buf_1
Xoutput42 net42 uo_out[7] VPWR VGND sg13g2_buf_1
Xheichips25_sap3__2782_ heichips25_sap3/_0427_ heichips25_sap3/_0425_ heichips25_sap3/_1605_
+ heichips25_sap3/_1762_ heichips25_sap3/_1643_ VPWR VGND sg13g2_a22oi_1
Xoutput31 net31 uio_out[4] VPWR VGND sg13g2_buf_1
Xoutput20 net20 uio_oe[1] VPWR VGND sg13g2_buf_1
Xheichips25_sap3_fanout95 heichips25_sap3/_1144_ heichips25_sap3/net95 VPWR VGND sg13g2_buf_1
Xheichips25_sap3_fanout73 heichips25_sap3/net74 heichips25_sap3/net73 VPWR VGND sg13g2_buf_1
XFILLER_1_742 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3403_ heichips25_sap3/_1010_ heichips25_sap3/net132 heichips25_sap3__3993_/Q
+ heichips25_sap3/net136 heichips25_sap3__3969_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_0_285 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3334_ heichips25_sap3/net52 heichips25_sap3/net50 heichips25_sap3/net48
+ heichips25_sap3/_0944_ VPWR VGND heichips25_sap3/_0943_ sg13g2_nand4_1
XFILLER_45_974 VPWR VGND sg13g2_decap_4
XFILLER_45_952 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3265_ heichips25_sap3/_1538_ heichips25_sap3/_0709_ heichips25_sap3/_0727_
+ heichips25_sap3/_0877_ heichips25_sap3/_0878_ VPWR VGND sg13g2_nor4_1
Xheichips25_sap3__3196_ heichips25_sap3/_0809_ heichips25_sap3/net104 heichips25_sap3__3951_/Q
+ heichips25_sap3/net144 heichips25_sap3__3967_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2216_ heichips25_sap3/_1636_ VPWR heichips25_sap3/_1637_ VGND heichips25_sap3/net236
+ heichips25_sap3/_1603_ sg13g2_o21ai_1
XFILLER_16_142 VPWR VGND sg13g2_fill_2
XFILLER_16_197 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2781__645 VPWR VGND net644 sg13g2_tiehi
Xheichips25_sap3__2147_ heichips25_sap3/_1547_ heichips25_sap3/_1567_ heichips25_sap3/_1568_
+ VPWR VGND sg13g2_nor2_1
XFILLER_31_145 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2078_ heichips25_sap3/_1499_ heichips25_sap3/net235 heichips25_sap3/net229
+ VPWR VGND sg13g2_nand2_1
XFILLER_12_381 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2933__604 VPWR VGND net603 sg13g2_tiehi
XFILLER_28_1028 VPWR VGND sg13g2_fill_1
XFILLER_39_212 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2822_ net562 VGND VPWR heichips25_can_lehmann_fsm/net1185
+ heichips25_can_lehmann_fsm__2822_/Q clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_39_267 VPWR VGND sg13g2_decap_8
XFILLER_39_278 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2753_ VGND VPWR heichips25_can_lehmann_fsm/_0856_ heichips25_can_lehmann_fsm/net386
+ heichips25_can_lehmann_fsm/_0276_ heichips25_can_lehmann_fsm/_0842_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2684_ heichips25_can_lehmann_fsm/net465 VPWR heichips25_can_lehmann_fsm/_0808_
+ VGND heichips25_can_lehmann_fsm__3016_/Q heichips25_can_lehmann_fsm/net358 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__1704_ heichips25_can_lehmann_fsm/_1028_ heichips25_can_lehmann_fsm/_1023_
+ heichips25_can_lehmann_fsm/_1027_ heichips25_can_lehmann_fsm/net300 heichips25_can_lehmann_fsm/_0953_
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2827__553 VPWR VGND net552 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__1635_ VPWR heichips25_can_lehmann_fsm/_0959_ heichips25_can_lehmann_fsm/net942
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__1566_ VPWR heichips25_can_lehmann_fsm/_0890_ heichips25_can_lehmann_fsm/net1021
+ VGND sg13g2_inv_1
XFILLER_10_329 VPWR VGND sg13g2_fill_1
XFILLER_31_690 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2118_ VGND VPWR heichips25_can_lehmann_fsm__2999_/Q heichips25_can_lehmann_fsm/net317
+ heichips25_can_lehmann_fsm/_0457_ heichips25_can_lehmann_fsm/net301 sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2049_ heichips25_can_lehmann_fsm/_1060_ heichips25_can_lehmann_fsm__2793_/Q
+ heichips25_can_lehmann_fsm/_0397_ VPWR VGND sg13g2_xor2_1
XFILLER_39_790 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3050_ VPWR heichips25_sap3/_0663_ heichips25_sap3/_0662_ VGND sg13g2_inv_1
XFILLER_13_101 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2001_ VPWR heichips25_sap3/_1427_ heichips25_sap3/net1128 VGND sg13g2_inv_1
XFILLER_41_443 VPWR VGND sg13g2_fill_1
XFILLER_13_167 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3952_ heichips25_sap3/net441 VGND VPWR heichips25_sap3/_0093_ heichips25_sap3__3952_/Q
+ clkload20/A sg13g2_dfrbpq_1
Xheichips25_sap3__2903_ VPWR VGND heichips25_sap3/net280 heichips25_sap3/_0542_ heichips25_sap3/_0417_
+ heichips25_sap3/net276 heichips25_sap3/_0543_ heichips25_sap3/_0416_ sg13g2_a221oi_1
XFILLER_6_867 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3883_ heichips25_sap3/net450 VGND VPWR heichips25_sap3/_0024_ heichips25_sap3__3883_/Q
+ heichips25_sap3__3922_/CLK sg13g2_dfrbpq_1
Xheichips25_sap3__2834_ heichips25_sap3/_0360_ heichips25_sap3/_0449_ heichips25_sap3/_0477_
+ VPWR VGND sg13g2_and2_1
Xheichips25_sap3__2765_ VGND VPWR heichips25_sap3/net276 heichips25_sap3/_1398_ heichips25_sap3/_0411_
+ heichips25_sap3/_0398_ sg13g2_a21oi_1
XFILLER_3_35 VPWR VGND sg13g2_decap_8
XFILLER_49_532 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2696_ heichips25_sap3/_0342_ heichips25_sap3/_0339_ heichips25_sap3/_0341_
+ VPWR VGND sg13g2_nand2_1
XFILLER_3_1019 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3317_ heichips25_sap3/_0928_ heichips25_sap3/_0909_ heichips25_sap3/net50
+ VPWR VGND sg13g2_xnor2_1
XFILLER_17_451 VPWR VGND sg13g2_fill_2
XFILLER_44_281 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3248_ heichips25_sap3/_0861_ heichips25_sap3/net122 heichips25_sap3/_0860_
+ VPWR VGND sg13g2_nand2_1
XFILLER_32_432 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3179_ heichips25_sap3/_0792_ heichips25_sap3__3969_/Q heichips25_sap3/net144
+ VPWR VGND sg13g2_nand2_1
XFILLER_33_988 VPWR VGND sg13g2_fill_1
XFILLER_32_498 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__3021_ net714 VGND VPWR heichips25_can_lehmann_fsm/_0246_
+ heichips25_can_lehmann_fsm__3021_/Q clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_41_1025 VPWR VGND sg13g2_decap_4
XFILLER_27_204 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2805_ net596 VGND VPWR heichips25_can_lehmann_fsm/net1203
+ heichips25_can_lehmann_fsm__2805_/Q clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_27_248 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2736_ heichips25_can_lehmann_fsm/net467 VPWR heichips25_can_lehmann_fsm/_0834_
+ VGND heichips25_can_lehmann_fsm__3043_/Q heichips25_can_lehmann_fsm/net391 sg13g2_o21ai_1
XFILLER_36_793 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2667_ VGND VPWR heichips25_can_lehmann_fsm/_0879_ heichips25_can_lehmann_fsm/net415
+ heichips25_can_lehmann_fsm/_0233_ heichips25_can_lehmann_fsm/_0799_ sg13g2_a21oi_1
XFILLER_10_115 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1618_ VPWR heichips25_can_lehmann_fsm/_0942_ heichips25_can_lehmann_fsm/net1177
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__2598_ heichips25_can_lehmann_fsm/net493 VPWR heichips25_can_lehmann_fsm/_0765_
+ VGND heichips25_can_lehmann_fsm__2974_/Q heichips25_can_lehmann_fsm/net407 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm_hold859 heichips25_can_lehmann_fsm__2929_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net858 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold848 heichips25_can_lehmann_fsm/_0201_ VPWR VGND heichips25_can_lehmann_fsm/net847
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__1549_ VPWR heichips25_can_lehmann_fsm/_0873_ heichips25_can_lehmann_fsm/net990
+ VGND sg13g2_inv_1
XFILLER_12_44 VPWR VGND sg13g2_fill_1
XFILLER_3_804 VPWR VGND sg13g2_decap_4
XFILLER_12_88 VPWR VGND sg13g2_decap_8
XFILLER_2_347 VPWR VGND sg13g2_decap_4
Xclkbuf_5_20__f_heichips25_sap3\_sap_3_inst.alu_inst.clk heichips25_sap3__3921_/CLK
+ clknet_4_10_0_heichips25_sap3\/sap_3_inst.alu_inst.clk VPWR VGND sg13g2_buf_16
Xheichips25_sap3__2550_ heichips25_sap3/_0225_ heichips25_sap3/net73 heichips25_sap3__3998_/Q
+ heichips25_sap3/net77 heichips25_sap3__4014_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2481_ heichips25_sap3/_1884_ heichips25_sap3/net168 heichips25_sap3/_1894_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__3102_ VGND VPWR heichips25_sap3/net247 heichips25_sap3/net246 heichips25_sap3/_0715_
+ heichips25_sap3/_0654_ sg13g2_a21oi_1
XFILLER_14_410 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3033_ heichips25_sap3/_0646_ heichips25_sap3/_1644_ heichips25_sap3/_1762_
+ VPWR VGND sg13g2_nand2_1
XFILLER_42_785 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3935_ heichips25_sap3/net438 VGND VPWR heichips25_sap3/_0076_ heichips25_sap3__3935_/Q
+ heichips25_sap3__4017_/CLK sg13g2_dfrbpq_1
Xheichips25_sap3__3866_ heichips25_sap3__3885_/Q heichips25_sap3/net1119 heichips25_sap3/net341
+ heichips25_sap3/_0193_ VPWR VGND sg13g2_mux2_1
Xheichips25_sap3__2817_ heichips25_sap3/_1381_ heichips25_sap3/_1619_ heichips25_sap3/_1714_
+ heichips25_sap3/_0461_ VPWR VGND sg13g2_nor3_1
XFILLER_5_196 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3797_ heichips25_sap3/_1306_ heichips25_sap3/_1279_ heichips25_sap3__3966_/Q
+ heichips25_sap3/net293 heichips25_sap3__3990_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2748_ VGND VPWR heichips25_sap3/_0387_ heichips25_sap3/_0393_ heichips25_sap3/_0394_
+ heichips25_sap3/_0388_ sg13g2_a21oi_1
Xheichips25_sap3__2679_ heichips25_sap3/_0330_ heichips25_sap3__3885_/Q heichips25_sap3/net213
+ VPWR VGND sg13g2_nand2_1
XFILLER_37_502 VPWR VGND sg13g2_fill_1
XFILLER_45_590 VPWR VGND sg13g2_decap_4
XFILLER_17_270 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2521_ VGND VPWR heichips25_can_lehmann_fsm/_0917_ heichips25_can_lehmann_fsm/net376
+ heichips25_can_lehmann_fsm/_0160_ heichips25_can_lehmann_fsm/_0726_ sg13g2_a21oi_1
XFILLER_32_240 VPWR VGND sg13g2_decap_8
XFILLER_21_925 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2452_ heichips25_can_lehmann_fsm/net472 VPWR heichips25_can_lehmann_fsm/_0692_
+ VGND heichips25_can_lehmann_fsm__2900_/Q heichips25_can_lehmann_fsm/net365 sg13g2_o21ai_1
XFILLER_32_251 VPWR VGND sg13g2_fill_1
XFILLER_21_958 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2383_ VGND VPWR heichips25_can_lehmann_fsm/_0956_ heichips25_can_lehmann_fsm/net423
+ heichips25_can_lehmann_fsm/_0091_ heichips25_can_lehmann_fsm/_0657_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm_fanout501 heichips25_can_lehmann_fsm/net502 heichips25_can_lehmann_fsm/net501
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm__3004_ net561 VGND VPWR heichips25_can_lehmann_fsm/_0229_
+ heichips25_can_lehmann_fsm__3004_/Q clknet_leaf_11_clk sg13g2_dfrbpq_1
Xclkbuf_4_5_0_heichips25_sap3\_sap_3_inst.alu_inst.clk clknet_0_heichips25_sap3\/sap_3_inst.alu_inst.clk
+ clknet_4_5_0_heichips25_sap3\/sap_3_inst.alu_inst.clk VPWR VGND sg13g2_buf_8
XFILLER_43_516 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2985__685 VPWR VGND net684 sg13g2_tiehi
XFILLER_28_568 VPWR VGND sg13g2_fill_1
XFILLER_43_549 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2719_ VGND VPWR heichips25_can_lehmann_fsm/_0865_ heichips25_can_lehmann_fsm/net371
+ heichips25_can_lehmann_fsm/_0259_ heichips25_can_lehmann_fsm/_0825_ sg13g2_a21oi_1
XFILLER_23_10 VPWR VGND sg13g2_fill_1
XFILLER_23_251 VPWR VGND sg13g2_fill_2
XFILLER_24_796 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__1981_ VPWR heichips25_sap3/_1407_ heichips25_sap3__4000_/Q VGND
+ sg13g2_inv_1
Xheichips25_sap3__3720_ heichips25_sap3__4021_/Q heichips25_sap3/_1066_ heichips25_sap3/net117
+ heichips25_sap3/_0162_ VPWR VGND sg13g2_mux2_1
XFILLER_2_111 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3651_ VGND VPWR heichips25_sap3/net48 heichips25_sap3/net51 heichips25_sap3/_1199_
+ heichips25_sap3/_0889_ sg13g2_a21oi_1
Xheichips25_sap3__2602_ heichips25_sap3__3901_/Q heichips25_sap3/net283 heichips25_sap3/_0274_
+ VPWR VGND sg13g2_xor2_1
Xheichips25_sap3__3582_ heichips25_sap3/_0107_ heichips25_sap3/_1107_ heichips25_sap3/_1158_
+ heichips25_sap3/net100 heichips25_sap3/_1372_ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2533_ heichips25_sap3/_1742_ heichips25_sap3/_0207_ heichips25_sap3/_0208_
+ heichips25_sap3/_0209_ heichips25_sap3/_0210_ VPWR VGND sg13g2_and4_1
Xheichips25_sap3__2464_ heichips25_sap3/_1877_ heichips25_sap3/_1873_ heichips25_sap3/_1876_
+ heichips25_sap3/_1869_ heichips25_sap3/_1866_ VPWR VGND sg13g2_a22oi_1
XFILLER_0_14 VPWR VGND sg13g2_fill_2
XFILLER_0_58 VPWR VGND sg13g2_decap_8
XFILLER_0_47 VPWR VGND sg13g2_fill_1
XFILLER_0_36 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2395_ heichips25_sap3/_1814_ heichips25_sap3__3896_/Q heichips25_sap3/_1788_
+ VPWR VGND sg13g2_nand2_1
XFILLER_34_549 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2964__769 VPWR VGND net768 sg13g2_tiehi
XFILLER_15_730 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__4065_ heichips25_sap3/net433 VGND VPWR heichips25_sap3/_0005_ heichips25_sap3__4065_/Q
+ net824 sg13g2_dfrbpq_1
XFILLER_9_45 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3016_ heichips25_sap3/_0634_ heichips25_sap3/net265 heichips25_sap3/net232
+ VPWR VGND sg13g2_nand2_1
XFILLER_30_744 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3918_ heichips25_sap3/net449 VGND VPWR heichips25_sap3/_0059_ heichips25_sap3__3918_/Q
+ heichips25_sap3__3920_/CLK sg13g2_dfrbpq_1
Xheichips25_sap3__3849_ heichips25_sap3__4047_/Q heichips25_sap3__4056_/Q heichips25_sap3/_1349_
+ VPWR VGND heichips25_sap3/net342 sg13g2_nand3b_1
Xheichips25_can_lehmann_fsm__1952_ heichips25_can_lehmann_fsm/net322 VPWR heichips25_can_lehmann_fsm/_0315_
+ VGND heichips25_can_lehmann_fsm/net1242 heichips25_can_lehmann_fsm/net179 sg13g2_o21ai_1
XFILLER_37_332 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1883_ VPWR VGND heichips25_can_lehmann_fsm/_1163_ heichips25_can_lehmann_fsm/_1195_
+ heichips25_can_lehmann_fsm/_1196_ heichips25_can_lehmann_fsm/net1164 heichips25_can_lehmann_fsm/_1197_
+ heichips25_can_lehmann_fsm/_1166_ sg13g2_a221oi_1
XFILLER_25_516 VPWR VGND sg13g2_decap_8
Xheichips25_sap3_fanout438 heichips25_sap3/net446 heichips25_sap3/net438 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout449 heichips25_sap3/net463 heichips25_sap3/net449 VPWR VGND
+ sg13g2_buf_1
Xheichips25_can_lehmann_fsm__2504_ heichips25_can_lehmann_fsm/net493 VPWR heichips25_can_lehmann_fsm/_0718_
+ VGND heichips25_can_lehmann_fsm/net1092 heichips25_can_lehmann_fsm/net366 sg13g2_o21ai_1
XFILLER_21_755 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__3002__578 VPWR VGND net577 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2435_ VGND VPWR heichips25_can_lehmann_fsm/_0939_ heichips25_can_lehmann_fsm/net409
+ heichips25_can_lehmann_fsm/_0117_ heichips25_can_lehmann_fsm/_0683_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2366_ heichips25_can_lehmann_fsm/net501 VPWR heichips25_can_lehmann_fsm/_0649_
+ VGND heichips25_can_lehmann_fsm/net968 heichips25_can_lehmann_fsm/net430 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2297_ heichips25_can_lehmann_fsm/_1051_ heichips25_can_lehmann_fsm/net209
+ heichips25_can_lehmann_fsm/_0608_ VPWR VGND sg13g2_nor2b_1
Xheichips25_can_lehmann_fsm_fanout320 heichips25_can_lehmann_fsm/_0990_ heichips25_can_lehmann_fsm/net320
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout331 heichips25_can_lehmann_fsm/net334 heichips25_can_lehmann_fsm/net331
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout364 heichips25_can_lehmann_fsm/net389 heichips25_can_lehmann_fsm/net364
+ VPWR VGND sg13g2_buf_1
XFILLER_0_604 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm_fanout375 heichips25_can_lehmann_fsm/net379 heichips25_can_lehmann_fsm/net375
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout353 heichips25_can_lehmann_fsm/net354 heichips25_can_lehmann_fsm/net353
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout386 heichips25_can_lehmann_fsm/net387 heichips25_can_lehmann_fsm/net386
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout397 heichips25_can_lehmann_fsm/net400 heichips25_can_lehmann_fsm/net397
+ VPWR VGND sg13g2_buf_1
XFILLER_28_332 VPWR VGND sg13g2_fill_2
XFILLER_18_76 VPWR VGND sg13g2_decap_8
XFILLER_43_335 VPWR VGND sg13g2_fill_1
XFILLER_43_324 VPWR VGND sg13g2_fill_1
XFILLER_43_302 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2180_ heichips25_sap3/net266 heichips25_sap3/_1510_ heichips25_sap3/_1553_
+ heichips25_sap3/_1601_ VPWR VGND sg13g2_nor3_1
XFILLER_43_346 VPWR VGND sg13g2_fill_2
XFILLER_31_508 VPWR VGND sg13g2_decap_4
XFILLER_24_560 VPWR VGND sg13g2_decap_8
XFILLER_8_704 VPWR VGND sg13g2_fill_2
XFILLER_12_744 VPWR VGND sg13g2_decap_4
XFILLER_15_1019 VPWR VGND sg13g2_fill_1
XFILLER_24_593 VPWR VGND sg13g2_fill_1
XFILLER_7_214 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__1964_ VPWR heichips25_sap3/_1390_ heichips25_sap3__3956_/Q VGND
+ sg13g2_inv_1
XFILLER_4_987 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2890__716 VPWR VGND net715 sg13g2_tiehi
Xheichips25_sap3__3703_ heichips25_sap3/_0153_ heichips25_sap3/_1095_ heichips25_sap3/_1234_
+ heichips25_sap3/net115 heichips25_sap3/_1386_ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3634_ heichips25_sap3/_1190_ heichips25_sap3__3988_/Q heichips25_sap3/net93
+ VPWR VGND sg13g2_nand2_1
XFILLER_38_118 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3565_ VGND VPWR heichips25_sap3/_0212_ heichips25_sap3/net95 heichips25_sap3/_1146_
+ heichips25_sap3/_1145_ sg13g2_a21oi_1
Xheichips25_sap3__2516_ heichips25_sap3/_1927_ heichips25_sap3/net71 heichips25_sap3__3971_/Q
+ heichips25_sap3/net216 heichips25_sap3__4003_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3496_ heichips25_sap3/_1084_ VPWR heichips25_sap3/_0088_ VGND heichips25_sap3/_1085_
+ heichips25_sap3/_1092_ sg13g2_o21ai_1
Xheichips25_sap3__2447_ heichips25_sap3/_1862_ heichips25_sap3/net77 heichips25_sap3__4023_/Q
+ heichips25_sap3/net84 heichips25_sap3__3967_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2929__620 VPWR VGND net619 sg13g2_tiehi
XFILLER_34_302 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2378_ heichips25_sap3/_1799_ heichips25_sap3/_1796_ heichips25_sap3/_1797_
+ heichips25_sap3/_1798_ VPWR VGND sg13g2_and3_1
XFILLER_22_519 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__4048_ heichips25_sap3/net452 VGND VPWR heichips25_sap3/_0189_ heichips25_sap3__4048_/Q
+ clknet_leaf_22_clk sg13g2_dfrbpq_1
XFILLER_30_574 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2220_ VGND VPWR heichips25_can_lehmann_fsm/net162 heichips25_can_lehmann_fsm/_0545_
+ heichips25_can_lehmann_fsm/_0039_ heichips25_can_lehmann_fsm/_0546_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2151_ heichips25_can_lehmann_fsm/_0490_ heichips25_can_lehmann_fsm__3046_/Q
+ heichips25_can_lehmann_fsm/_1161_ VPWR VGND sg13g2_nand2_1
Xheichips25_can_lehmann_fsm__2082_ VPWR VGND heichips25_can_lehmann_fsm/_0425_ heichips25_can_lehmann_fsm/_1176_
+ heichips25_can_lehmann_fsm/_0424_ heichips25_can_lehmann_fsm/_0976_ heichips25_can_lehmann_fsm/_0022_
+ heichips25_can_lehmann_fsm/net182 sg13g2_a221oi_1
Xheichips25_can_lehmann_fsm__2791__625 VPWR VGND net624 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__3010__803 VPWR VGND net802 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2984_ net688 VGND VPWR heichips25_can_lehmann_fsm/_0209_
+ heichips25_can_lehmann_fsm__2984_/Q clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_29_129 VPWR VGND sg13g2_fill_2
XFILLER_37_140 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1935_ heichips25_can_lehmann_fsm/_0298_ heichips25_can_lehmann_fsm/net312
+ heichips25_can_lehmann_fsm__3026_/Q heichips25_can_lehmann_fsm/net319 heichips25_can_lehmann_fsm__3002_/Q
+ VPWR VGND sg13g2_a22oi_1
XFILLER_37_173 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1866_ heichips25_can_lehmann_fsm/_1181_ heichips25_can_lehmann_fsm/net297
+ heichips25_can_lehmann_fsm__2891_/Q heichips25_can_lehmann_fsm/net314 heichips25_can_lehmann_fsm__2915_/Q
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3_fanout213 heichips25_sap3/net214 heichips25_sap3/net213 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout202 heichips25_sap3/_0624_ heichips25_sap3/net202 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout235 heichips25_sap3/_1462_ heichips25_sap3/net235 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout224 heichips25_sap3/_1622_ heichips25_sap3/net224 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout257 heichips25_sap3/_1362_ heichips25_sap3/net257 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout246 heichips25_sap3/_1467_ heichips25_sap3/net246 VPWR VGND
+ sg13g2_buf_1
XFILLER_25_335 VPWR VGND sg13g2_fill_1
Xheichips25_sap3_fanout268 heichips25_sap3__3925_/Q heichips25_sap3/net268 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout279 heichips25_sap3__3904_/Q heichips25_sap3/net279 VPWR VGND
+ sg13g2_buf_1
Xheichips25_can_lehmann_fsm__1797_ VPWR VGND heichips25_can_lehmann_fsm__2901_/Q heichips25_can_lehmann_fsm/_1112_
+ heichips25_can_lehmann_fsm/net296 heichips25_can_lehmann_fsm__2925_/Q heichips25_can_lehmann_fsm/_1113_
+ heichips25_can_lehmann_fsm/net313 sg13g2_a221oi_1
Xheichips25_can_lehmann_fsm__2418_ heichips25_can_lehmann_fsm/net497 VPWR heichips25_can_lehmann_fsm/_0675_
+ VGND heichips25_can_lehmann_fsm/net977 heichips25_can_lehmann_fsm/net384 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2349_ VGND VPWR heichips25_can_lehmann_fsm/_0964_ heichips25_can_lehmann_fsm/net382
+ heichips25_can_lehmann_fsm/_0074_ heichips25_can_lehmann_fsm/_0640_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2837__533 VPWR VGND net532 sg13g2_tiehi
Xheichips25_can_lehmann_fsm_fanout172 heichips25_can_lehmann_fsm/net173 heichips25_can_lehmann_fsm/net172
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout161 heichips25_can_lehmann_fsm/net163 heichips25_can_lehmann_fsm/net161
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout183 heichips25_can_lehmann_fsm/_0312_ heichips25_can_lehmann_fsm/net183
+ VPWR VGND sg13g2_buf_1
XFILLER_20_88 VPWR VGND sg13g2_fill_2
XFILLER_1_968 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm_fanout194 heichips25_can_lehmann_fsm/_0306_ heichips25_can_lehmann_fsm/net194
+ VPWR VGND sg13g2_buf_1
Xheichips25_sap3__3350_ VPWR VGND heichips25_sap3__3999_/Q heichips25_sap3/net129
+ heichips25_sap3/net148 heichips25_sap3__4015_/Q heichips25_sap3/_0959_ heichips25_sap3/net116
+ sg13g2_a221oi_1
XFILLER_29_86 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2301_ heichips25_sap3/_1722_ heichips25_sap3/net264 heichips25_sap3/net256
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__3281_ heichips25_sap3/_0893_ heichips25_sap3/net145 heichips25_sap3__3956_/Q
+ heichips25_sap3/net146 heichips25_sap3__3996_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2232_ heichips25_sap3/_1653_ heichips25_sap3/_1471_ heichips25_sap3/_1652_
+ VPWR VGND sg13g2_nand2_1
XFILLER_28_184 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__3022__707 VPWR VGND net706 sg13g2_tiehi
Xheichips25_sap3__2163_ heichips25_sap3/_1584_ heichips25_sap3/_1582_ heichips25_sap3/_1575_
+ VPWR VGND sg13g2_nand2b_1
Xheichips25_sap3__2094_ heichips25_sap3/net261 heichips25_sap3/_1446_ heichips25_sap3/_1506_
+ heichips25_sap3/_1515_ VPWR VGND sg13g2_nor3_1
XFILLER_31_338 VPWR VGND sg13g2_decap_8
XFILLER_31_349 VPWR VGND sg13g2_fill_1
XFILLER_12_541 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3880__825 VPWR net824 heichips25_sap3__4013_/CLK VGND sg13g2_inv_1
Xheichips25_sap3__2996_ heichips25_sap3__3915_/Q heichips25_sap3/net201 heichips25_sap3/_0625_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__1947_ VPWR heichips25_sap3/_1373_ heichips25_sap3__3950_/Q VGND
+ sg13g2_inv_1
XFILLER_3_294 VPWR VGND sg13g2_fill_1
XFILLER_6_1028 VPWR VGND sg13g2_fill_1
XFILLER_6_1006 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3617_ VGND VPWR heichips25_sap3/_1388_ heichips25_sap3/net102 heichips25_sap3/_0121_
+ heichips25_sap3/_1180_ sg13g2_a21oi_1
Xheichips25_sap3__3548_ heichips25_sap3/net56 VPWR heichips25_sap3/_1136_ VGND heichips25_sap3/_1061_
+ heichips25_sap3/_1062_ sg13g2_o21ai_1
Xheichips25_sap3__3479_ VGND VPWR heichips25_sap3/_1078_ heichips25_sap3/_1076_ net43
+ sg13g2_or2_1
XFILLER_19_162 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1720_ heichips25_can_lehmann_fsm/_1042_ heichips25_can_lehmann_fsm/_1037_
+ heichips25_can_lehmann_fsm__2787_/Q heichips25_can_lehmann_fsm/_1032_ heichips25_can_lehmann_fsm/net346
+ VPWR VGND sg13g2_a22oi_1
XFILLER_34_110 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__1651_ VPWR heichips25_can_lehmann_fsm/_0975_ heichips25_can_lehmann_fsm/net1226
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__1582_ VPWR heichips25_can_lehmann_fsm/_0906_ heichips25_can_lehmann_fsm/net1035
+ VGND sg13g2_inv_1
XFILLER_31_861 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2203_ VGND VPWR heichips25_can_lehmann_fsm/net163 heichips25_can_lehmann_fsm/_0532_
+ heichips25_can_lehmann_fsm/_0035_ heichips25_can_lehmann_fsm/_0533_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2134_ VPWR VGND heichips25_can_lehmann_fsm__2910_/Q heichips25_can_lehmann_fsm/_0472_
+ heichips25_can_lehmann_fsm/net298 heichips25_can_lehmann_fsm__3030_/Q heichips25_can_lehmann_fsm/_0473_
+ heichips25_can_lehmann_fsm/net312 sg13g2_a221oi_1
Xheichips25_can_lehmann_fsm__2065_ heichips25_can_lehmann_fsm/_0412_ heichips25_can_lehmann_fsm/_0411_
+ heichips25_can_lehmann_fsm/net189 VPWR VGND sg13g2_nand2b_1
XFILLER_39_983 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2967_ net756 VGND VPWR heichips25_can_lehmann_fsm/net886
+ heichips25_can_lehmann_fsm__2967_/Q clknet_leaf_20_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2898_ net699 VGND VPWR heichips25_can_lehmann_fsm/net914
+ heichips25_can_lehmann_fsm__2898_/Q clknet_leaf_21_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1918_ heichips25_can_lehmann_fsm/_1230_ VPWR heichips25_can_lehmann_fsm/_1231_
+ VGND heichips25_can_lehmann_fsm__2883_/Q heichips25_can_lehmann_fsm/net335 sg13g2_o21ai_1
XFILLER_13_305 VPWR VGND sg13g2_fill_2
XFILLER_15_22 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1849_ heichips25_can_lehmann_fsm/_1090_ VPWR heichips25_can_lehmann_fsm/_1165_
+ VGND heichips25_can_lehmann_fsm/_1096_ heichips25_can_lehmann_fsm/_1164_ sg13g2_o21ai_1
XFILLER_25_154 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm_hold1100 heichips25_can_lehmann_fsm__2839_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1099 sg13g2_dlygate4sd3_1
XFILLER_40_135 VPWR VGND sg13g2_decap_8
XFILLER_15_33 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_hold1133 heichips25_can_lehmann_fsm__3059_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1132 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1111 heichips25_can_lehmann_fsm__2876_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1110 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1166 heichips25_can_lehmann_fsm__2829_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1165 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1155 heichips25_can_lehmann_fsm__3045_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1154 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1188 heichips25_can_lehmann_fsm/_0038_ VPWR VGND heichips25_can_lehmann_fsm/net1187
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1199 heichips25_can_lehmann_fsm__2809_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1198 sg13g2_dlygate4sd3_1
Xheichips25_sap3_hold831 heichips25_sap3__4059_/Q VPWR VGND heichips25_sap3/net830
+ sg13g2_dlygate4sd3_1
XFILLER_31_43 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2850_ heichips25_sap3/net64 heichips25_sap3/_0477_ heichips25_sap3/_0479_
+ heichips25_sap3/_0492_ heichips25_sap3/_0493_ VPWR VGND sg13g2_or4_1
Xheichips25_sap3_fanout63 heichips25_sap3/_0810_ heichips25_sap3/net63 VPWR VGND sg13g2_buf_1
Xheichips25_sap3_fanout52 heichips25_sap3/_0898_ heichips25_sap3/net52 VPWR VGND sg13g2_buf_1
Xheichips25_sap3_fanout96 heichips25_sap3/net97 heichips25_sap3/net96 VPWR VGND sg13g2_buf_1
Xheichips25_sap3__2781_ heichips25_sap3/net223 heichips25_sap3/_1727_ heichips25_sap3/_0426_
+ VPWR VGND sg13g2_nor2_1
Xoutput32 net32 uio_out[5] VPWR VGND sg13g2_buf_1
Xoutput21 net21 uio_oe[2] VPWR VGND sg13g2_buf_1
Xheichips25_sap3_fanout74 heichips25_sap3/_1745_ heichips25_sap3/net74 VPWR VGND sg13g2_buf_2
Xheichips25_sap3_fanout85 heichips25_sap3/net86 heichips25_sap3/net85 VPWR VGND sg13g2_buf_1
XFILLER_0_220 VPWR VGND sg13g2_decap_8
XFILLER_0_253 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3402_ heichips25_sap3/_1009_ heichips25_sap3__3945_/Q heichips25_sap3/_0763_
+ VPWR VGND sg13g2_nand2_1
XFILLER_0_297 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3333_ VGND VPWR heichips25_sap3/_1368_ heichips25_sap3/net127 heichips25_sap3/_0943_
+ heichips25_sap3/_0942_ sg13g2_a21oi_1
XFILLER_29_471 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3264_ heichips25_sap3/_1573_ VPWR heichips25_sap3/_0877_ VGND heichips25_sap3/_1527_
+ heichips25_sap3/_1569_ sg13g2_o21ai_1
Xheichips25_sap3__3195_ heichips25_sap3/_0808_ heichips25_sap3/net109 heichips25_sap3__3959_/Q
+ heichips25_sap3/net129 heichips25_sap3__3943_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2215_ heichips25_sap3/_1531_ heichips25_sap3/_1635_ heichips25_sap3/_1636_
+ VPWR VGND sg13g2_and2_1
XFILLER_17_677 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2146_ VGND VPWR heichips25_sap3/_1567_ heichips25_sap3/net252 heichips25_sap3/net253
+ sg13g2_or2_1
Xheichips25_sap3__2077_ heichips25_sap3/net236 heichips25_sap3/_1496_ heichips25_sap3/_1498_
+ VPWR VGND sg13g2_nor2_1
XFILLER_8_386 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2979_ heichips25_sap3/_0050_ heichips25_sap3/_0612_ heichips25_sap3/_0613_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_can_lehmann_fsm__2821_ net564 VGND VPWR heichips25_can_lehmann_fsm/_0046_
+ heichips25_can_lehmann_fsm__2821_/Q clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_39_246 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2752_ heichips25_can_lehmann_fsm/net499 VPWR heichips25_can_lehmann_fsm/_0842_
+ VGND heichips25_can_lehmann_fsm/net1157 heichips25_can_lehmann_fsm/net386 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__1703_ VPWR VGND heichips25_can_lehmann_fsm__2943_/Q heichips25_can_lehmann_fsm/_1026_
+ heichips25_can_lehmann_fsm/net305 heichips25_can_lehmann_fsm__3015_/Q heichips25_can_lehmann_fsm/_1027_
+ heichips25_can_lehmann_fsm/net310 sg13g2_a221oi_1
Xheichips25_can_lehmann_fsm__2683_ VGND VPWR heichips25_can_lehmann_fsm/_0875_ heichips25_can_lehmann_fsm/net397
+ heichips25_can_lehmann_fsm/_0241_ heichips25_can_lehmann_fsm/_0807_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__1634_ VPWR heichips25_can_lehmann_fsm/_0958_ heichips25_can_lehmann_fsm/net948
+ VGND sg13g2_inv_1
XFILLER_22_102 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__1565_ VPWR heichips25_can_lehmann_fsm/_0889_ heichips25_can_lehmann_fsm/net918
+ VGND sg13g2_inv_1
XFILLER_2_507 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2117_ heichips25_can_lehmann_fsm/_0456_ heichips25_can_lehmann_fsm/net294
+ heichips25_can_lehmann_fsm__2975_/Q heichips25_can_lehmann_fsm/net299 heichips25_can_lehmann_fsm__2903_/Q
+ VPWR VGND sg13g2_a22oi_1
XFILLER_7_9 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2048_ VGND VPWR heichips25_can_lehmann_fsm/net177 heichips25_can_lehmann_fsm/_0395_
+ heichips25_can_lehmann_fsm/_0017_ heichips25_can_lehmann_fsm/_0396_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__3051__799 VPWR VGND net798 sg13g2_tiehi
XFILLER_19_909 VPWR VGND sg13g2_decap_4
XFILLER_45_216 VPWR VGND sg13g2_fill_1
XFILLER_26_32 VPWR VGND sg13g2_fill_1
XFILLER_26_43 VPWR VGND sg13g2_fill_1
XFILLER_26_65 VPWR VGND sg13g2_decap_4
XFILLER_42_945 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2000_ VPWR heichips25_sap3/_1426_ heichips25_sap3__4038_/Q VGND
+ sg13g2_inv_1
XFILLER_26_485 VPWR VGND sg13g2_decap_8
XFILLER_14_669 VPWR VGND sg13g2_decap_8
XFILLER_42_53 VPWR VGND sg13g2_fill_1
XFILLER_41_488 VPWR VGND sg13g2_fill_1
XFILLER_41_477 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3951_ heichips25_sap3/net439 VGND VPWR heichips25_sap3/_0092_ heichips25_sap3__3951_/Q
+ clkload18/A sg13g2_dfrbpq_1
Xheichips25_sap3__2902_ heichips25_sap3/net278 heichips25_sap3/_0441_ heichips25_sap3/_0542_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_can_lehmann_fsm__3056__622 VPWR VGND net621 sg13g2_tiehi
Xheichips25_sap3__3882_ heichips25_sap3/net450 VGND VPWR heichips25_sap3/_0023_ heichips25_sap3__3882_/Q
+ heichips25_sap3__3922_/CLK sg13g2_dfrbpq_1
Xheichips25_sap3__2833_ net44 heichips25_sap3/net158 heichips25_sap3/_0476_ VPWR VGND
+ sg13g2_nor2b_1
Xheichips25_sap3__2764_ heichips25_sap3/_0399_ heichips25_sap3/_0409_ heichips25_sap3/_0410_
+ VPWR VGND sg13g2_nor2_1
XFILLER_1_540 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2695_ heichips25_sap3/_0341_ heichips25_sap3/_1886_ heichips25_sap3/_1892_
+ VPWR VGND sg13g2_nand2_1
XFILLER_3_58 VPWR VGND sg13g2_decap_8
XFILLER_49_555 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3316_ heichips25_sap3/net51 heichips25_sap3/net50 heichips25_sap3/net48
+ heichips25_sap3/_0927_ VPWR VGND sg13g2_nand3_1
Xheichips25_sap3__3247_ heichips25_sap3/_0860_ heichips25_sap3/_0777_ heichips25_sap3/_0858_
+ VPWR VGND sg13g2_xnor2_1
XFILLER_45_794 VPWR VGND sg13g2_fill_1
XFILLER_44_260 VPWR VGND sg13g2_fill_1
XFILLER_17_485 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3178_ heichips25_sap3/_0791_ heichips25_sap3__3953_/Q heichips25_sap3/net104
+ VPWR VGND sg13g2_nand2_1
XFILLER_33_978 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2129_ heichips25_sap3/_1550_ heichips25_sap3/net246 heichips25_sap3/_1546_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_can_lehmann_fsm__3020_ net722 VGND VPWR heichips25_can_lehmann_fsm/_0245_
+ heichips25_can_lehmann_fsm__3020_/Q clknet_leaf_0_clk sg13g2_dfrbpq_1
Xclkbuf_5_3__f_heichips25_sap3\_sap_3_inst.alu_inst.clk clkload18/A clknet_4_1_0_heichips25_sap3\/sap_3_inst.alu_inst.clk
+ VPWR VGND sg13g2_buf_16
Xheichips25_can_lehmann_fsm__2804_ net598 VGND VPWR heichips25_can_lehmann_fsm/net1216
+ heichips25_can_lehmann_fsm__2804_/Q clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_36_761 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2735_ VGND VPWR heichips25_can_lehmann_fsm/_0861_ heichips25_can_lehmann_fsm/net356
+ heichips25_can_lehmann_fsm/_0267_ heichips25_can_lehmann_fsm/_0833_ sg13g2_a21oi_1
XFILLER_35_271 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2666_ heichips25_can_lehmann_fsm/net483 VPWR heichips25_can_lehmann_fsm/_0799_
+ VGND heichips25_can_lehmann_fsm/net1150 heichips25_can_lehmann_fsm/net415 sg13g2_o21ai_1
XFILLER_23_433 VPWR VGND sg13g2_fill_1
XFILLER_23_466 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__3005__554 VPWR VGND net553 sg13g2_tiehi
Xheichips25_can_lehmann_fsm_hold849 heichips25_can_lehmann_fsm__3037_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net848 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__1617_ VPWR heichips25_can_lehmann_fsm/_0941_ heichips25_can_lehmann_fsm/net1003
+ VGND sg13g2_inv_1
XFILLER_23_499 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2597_ VGND VPWR heichips25_can_lehmann_fsm/_0898_ heichips25_can_lehmann_fsm/net366
+ heichips25_can_lehmann_fsm/_0198_ heichips25_can_lehmann_fsm/_0764_ sg13g2_a21oi_1
XFILLER_10_138 VPWR VGND sg13g2_decap_4
XFILLER_10_149 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1548_ VPWR heichips25_can_lehmann_fsm/_0872_ heichips25_can_lehmann_fsm/net1146
+ VGND sg13g2_inv_1
Xheichips25_sap3__2480_ heichips25_sap3/_1893_ heichips25_sap3/net168 heichips25_sap3/_1884_
+ VPWR VGND sg13g2_nand2b_1
XFILLER_18_205 VPWR VGND sg13g2_fill_1
XFILLER_37_64 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3101_ heichips25_sap3/_0314_ VPWR heichips25_sap3/_0714_ VGND heichips25_sap3/_1719_
+ heichips25_sap3/_0713_ sg13g2_o21ai_1
Xheichips25_sap3__3032_ heichips25_sap3/_1475_ heichips25_sap3/net226 heichips25_sap3/_1643_
+ heichips25_sap3/_0645_ VPWR VGND sg13g2_nor3_1
XFILLER_14_466 VPWR VGND sg13g2_fill_1
XFILLER_30_926 VPWR VGND sg13g2_fill_1
XFILLER_41_296 VPWR VGND sg13g2_decap_8
XFILLER_41_285 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3934_ heichips25_sap3/net438 VGND VPWR heichips25_sap3/_0075_ heichips25_sap3__3934_/Q
+ heichips25_sap3__4014_/CLK sg13g2_dfrbpq_1
Xheichips25_sap3__3865_ heichips25_sap3__3884_/Q heichips25_sap3/net1149 heichips25_sap3/net341
+ heichips25_sap3/_0192_ VPWR VGND sg13g2_mux2_1
XFILLER_5_175 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2816_ VGND VPWR heichips25_sap3/net154 heichips25_sap3/_0400_ heichips25_sap3/_0460_
+ heichips25_sap3/_0459_ sg13g2_a21oi_1
Xheichips25_sap3__3796_ VGND VPWR heichips25_sap3__3974_/Q heichips25_sap3/_1272_
+ heichips25_sap3/_1305_ heichips25_sap3/net290 sg13g2_a21oi_1
Xheichips25_sap3__2747_ VGND VPWR heichips25_sap3/net284 heichips25_sap3/_1397_ heichips25_sap3/_0393_
+ heichips25_sap3/_0392_ sg13g2_a21oi_1
Xheichips25_sap3__2678_ heichips25_sap3/net285 heichips25_sap3__3884_/Q heichips25_sap3/_0297_
+ heichips25_sap3/_0025_ VPWR VGND sg13g2_mux2_1
XFILLER_24_208 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2520_ heichips25_can_lehmann_fsm/net487 VPWR heichips25_can_lehmann_fsm/_0726_
+ VGND heichips25_can_lehmann_fsm__2934_/Q heichips25_can_lehmann_fsm/net378 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__3041__743 VPWR VGND net742 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2451_ VGND VPWR heichips25_can_lehmann_fsm/_0935_ heichips25_can_lehmann_fsm/net398
+ heichips25_can_lehmann_fsm/_0125_ heichips25_can_lehmann_fsm/_0691_ sg13g2_a21oi_1
XFILLER_32_263 VPWR VGND sg13g2_fill_1
XFILLER_33_786 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2382_ heichips25_can_lehmann_fsm/net495 VPWR heichips25_can_lehmann_fsm/_0657_
+ VGND heichips25_can_lehmann_fsm/net912 heichips25_can_lehmann_fsm/net423 sg13g2_o21ai_1
XFILLER_20_436 VPWR VGND sg13g2_fill_1
XFILLER_32_296 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm_fanout502 heichips25_can_lehmann_fsm/net503 heichips25_can_lehmann_fsm/net502
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm__3003_ net569 VGND VPWR heichips25_can_lehmann_fsm/net907
+ heichips25_can_lehmann_fsm__3003_/Q clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_28_503 VPWR VGND sg13g2_fill_1
XFILLER_28_547 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2718_ heichips25_can_lehmann_fsm/net478 VPWR heichips25_can_lehmann_fsm/_0825_
+ VGND heichips25_can_lehmann_fsm__3033_/Q heichips25_can_lehmann_fsm/net371 sg13g2_o21ai_1
XFILLER_24_753 VPWR VGND sg13g2_fill_2
XFILLER_23_274 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2649_ VGND VPWR heichips25_can_lehmann_fsm/_0884_ heichips25_can_lehmann_fsm/net404
+ heichips25_can_lehmann_fsm/_0224_ heichips25_can_lehmann_fsm/_0790_ sg13g2_a21oi_1
Xheichips25_sap3__1980_ VPWR heichips25_sap3/_1406_ heichips25_sap3__4008_/Q VGND
+ sg13g2_inv_1
Xheichips25_can_lehmann_fsm__2992__657 VPWR VGND net656 sg13g2_tiehi
Xheichips25_sap3__3650_ heichips25_sap3/net112 heichips25_sap3__3995_/Q heichips25_sap3/_1198_
+ heichips25_sap3/_0136_ VPWR VGND sg13g2_a21o_1
Xheichips25_sap3__2601_ heichips25_sap3/net289 heichips25_sap3/net287 heichips25_sap3/_0273_
+ VPWR VGND sg13g2_xor2_1
Xheichips25_sap3__3581_ heichips25_sap3/_1159_ heichips25_sap3/_0819_ heichips25_sap3/_0864_
+ VPWR VGND sg13g2_xnor2_1
Xheichips25_sap3__2532_ heichips25_sap3/_0209_ heichips25_sap3/net71 heichips25_sap3__3979_/Q
+ heichips25_sap3/net216 heichips25_sap3__4011_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_47_823 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2463_ heichips25_sap3/net221 heichips25_sap3/_1875_ heichips25_sap3/_1876_
+ VPWR VGND sg13g2_nor2_1
XFILLER_19_514 VPWR VGND sg13g2_fill_1
XFILLER_46_322 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2394_ heichips25_sap3/_1813_ net9 heichips25_sap3/_1770_ VPWR VGND
+ sg13g2_nand2_1
XFILLER_46_377 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__4064_ heichips25_sap3/net434 VGND VPWR heichips25_sap3/_0004_ heichips25_sap3__4064_/Q
+ net823 sg13g2_dfrbpq_1
Xheichips25_sap3__3015_ VGND VPWR heichips25_sap3/_1362_ heichips25_sap3/net231 heichips25_sap3/_0066_
+ heichips25_sap3/_0633_ sg13g2_a21oi_1
XFILLER_14_252 VPWR VGND sg13g2_decap_8
XFILLER_14_263 VPWR VGND sg13g2_fill_2
XFILLER_9_57 VPWR VGND sg13g2_fill_1
XFILLER_30_789 VPWR VGND sg13g2_fill_2
XFILLER_10_480 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3917_ heichips25_sap3/net447 VGND VPWR heichips25_sap3/_0058_ heichips25_sap3__3917_/Q
+ clkload24/A sg13g2_dfrbpq_1
XFILLER_43_4 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3848_ heichips25_sap3/net342 heichips25_sap3__4050_/Q heichips25_sap3__4051_/Q
+ heichips25_sap3__4052_/Q heichips25_sap3__4053_/Q heichips25_sap3__4047_/Q heichips25_sap3/_1348_
+ VPWR VGND sg13g2_mux4_1
Xheichips25_sap3__3779_ heichips25_sap3/_1290_ heichips25_sap3/net292 heichips25_sap3__3956_/Q
+ heichips25_sap3/net293 heichips25_sap3__3988_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__1951_ heichips25_can_lehmann_fsm/net347 heichips25_can_lehmann_fsm/net182
+ heichips25_can_lehmann_fsm/_0314_ VPWR VGND sg13g2_nor2_1
Xheichips25_can_lehmann_fsm__1882_ heichips25_can_lehmann_fsm/_1196_ heichips25_can_lehmann_fsm/_1153_
+ heichips25_can_lehmann_fsm/net305 VPWR VGND sg13g2_nand2b_1
Xheichips25_sap3_fanout439 heichips25_sap3/net446 heichips25_sap3/net439 VPWR VGND
+ sg13g2_buf_1
XFILLER_40_509 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2503_ VGND VPWR heichips25_can_lehmann_fsm/_0922_ heichips25_can_lehmann_fsm/net407
+ heichips25_can_lehmann_fsm/_0151_ heichips25_can_lehmann_fsm/_0717_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2434_ heichips25_can_lehmann_fsm/net477 VPWR heichips25_can_lehmann_fsm/_0683_
+ VGND heichips25_can_lehmann_fsm/net989 heichips25_can_lehmann_fsm/net410 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2365_ VGND VPWR heichips25_can_lehmann_fsm/_0960_ heichips25_can_lehmann_fsm/net387
+ heichips25_can_lehmann_fsm/_0082_ heichips25_can_lehmann_fsm/_0648_ sg13g2_a21oi_1
XFILLER_20_299 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2296_ heichips25_can_lehmann_fsm/_0607_ heichips25_can_lehmann_fsm/net206
+ heichips25_can_lehmann_fsm/net174 VPWR VGND sg13g2_nand2_1
Xheichips25_can_lehmann_fsm_fanout332 heichips25_can_lehmann_fsm/net334 heichips25_can_lehmann_fsm/net332
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout310 heichips25_can_lehmann_fsm/net312 heichips25_can_lehmann_fsm/net310
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout321 heichips25_can_lehmann_fsm/net324 heichips25_can_lehmann_fsm/net321
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout354 heichips25_can_lehmann_fsm__2775_/Q heichips25_can_lehmann_fsm/net354
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout343 heichips25_can_lehmann_fsm__3043_/Q heichips25_can_lehmann_fsm/net343
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout365 heichips25_can_lehmann_fsm/net367 heichips25_can_lehmann_fsm/net365
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout376 heichips25_can_lehmann_fsm/net379 heichips25_can_lehmann_fsm/net376
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout398 heichips25_can_lehmann_fsm/net399 heichips25_can_lehmann_fsm/net398
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout387 heichips25_can_lehmann_fsm/net388 heichips25_can_lehmann_fsm/net387
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm__2848__800 VPWR VGND net799 sg13g2_tiehi
XFILLER_28_355 VPWR VGND sg13g2_decap_8
XFILLER_34_43 VPWR VGND sg13g2_decap_8
XFILLER_11_222 VPWR VGND sg13g2_fill_2
XFILLER_34_87 VPWR VGND sg13g2_decap_8
XFILLER_34_98 VPWR VGND sg13g2_decap_8
XFILLER_11_255 VPWR VGND sg13g2_fill_2
XFILLER_7_226 VPWR VGND sg13g2_decap_8
Xclkbuf_5_21__f_heichips25_sap3\_sap_3_inst.alu_inst.clk clkload25/A clknet_4_10_0_heichips25_sap3\/sap_3_inst.alu_inst.clk
+ VPWR VGND sg13g2_buf_16
Xheichips25_sap3__1963_ VPWR heichips25_sap3/_1389_ heichips25_sap3__3964_/Q VGND
+ sg13g2_inv_1
Xheichips25_sap3__3702_ uio_oe_sap3\[1\] heichips25_sap3/net115 heichips25_sap3/_1234_
+ VPWR VGND sg13g2_nor2_1
XFILLER_1_0 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3633_ VPWR heichips25_sap3/_0128_ heichips25_sap3/_1189_ VGND sg13g2_inv_1
Xheichips25_sap3__3564_ uio_oe_sap3\[0\] heichips25_sap3/net95 heichips25_sap3/_1145_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__2515_ heichips25_sap3/_1926_ heichips25_sap3/net79 heichips25_sap3__4019_/Q
+ heichips25_sap3/net86 heichips25_sap3__3947_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3495_ heichips25_sap3/_1055_ heichips25_sap3/_1086_ heichips25_sap3/_1090_
+ heichips25_sap3/_1091_ heichips25_sap3/_1092_ VPWR VGND sg13g2_nor4_1
Xheichips25_sap3__2446_ heichips25_sap3/_1861_ heichips25_sap3/net85 heichips25_sap3__3959_/Q
+ heichips25_sap3/net87 heichips25_sap3__3951_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_46_185 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2377_ heichips25_sap3/_1798_ heichips25_sap3/net77 heichips25_sap3__4026_/Q
+ heichips25_sap3/net87 heichips25_sap3__3954_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__4047_ heichips25_sap3/net452 VGND VPWR heichips25_sap3/net1073 heichips25_sap3__4047_/Q
+ clknet_leaf_22_clk sg13g2_dfrbpq_1
XFILLER_15_583 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2150_ heichips25_can_lehmann_fsm/_1090_ VPWR heichips25_can_lehmann_fsm/_0489_
+ VGND heichips25_can_lehmann_fsm/_1138_ heichips25_can_lehmann_fsm/_0488_ sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2081_ heichips25_can_lehmann_fsm/_0425_ heichips25_can_lehmann_fsm/net195
+ net14 heichips25_can_lehmann_fsm/net199 heichips25_can_lehmann_fsm/net1219 VPWR
+ VGND sg13g2_a22oi_1
XFILLER_6_292 VPWR VGND sg13g2_fill_2
XFILLER_6_281 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2983_ net692 VGND VPWR heichips25_can_lehmann_fsm/net986
+ heichips25_can_lehmann_fsm__2983_/Q clknet_leaf_14_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1934_ heichips25_can_lehmann_fsm/_0297_ heichips25_can_lehmann_fsm/net333
+ heichips25_can_lehmann_fsm__3050_/Q heichips25_can_lehmann_fsm/net315 heichips25_can_lehmann_fsm__2930_/Q
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__1865_ heichips25_can_lehmann_fsm/_1180_ heichips25_can_lehmann_fsm/net295
+ heichips25_can_lehmann_fsm__2963_/Q heichips25_can_lehmann_fsm/net311 heichips25_can_lehmann_fsm__3011_/Q
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3_fanout214 heichips25_sap3/_0309_ heichips25_sap3/net214 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout203 heichips25_sap3/net204 heichips25_sap3/net203 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout236 heichips25_sap3/net240 heichips25_sap3/net236 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout225 heichips25_sap3/_1598_ heichips25_sap3/net225 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout247 heichips25_sap3/_1457_ heichips25_sap3/net247 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout258 heichips25_sap3__3930_/Q heichips25_sap3/net258 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout269 heichips25_sap3/net270 heichips25_sap3/net269 VPWR VGND
+ sg13g2_buf_1
Xheichips25_can_lehmann_fsm__1796_ heichips25_can_lehmann_fsm/net336 VPWR heichips25_can_lehmann_fsm/_1112_
+ VGND heichips25_can_lehmann_fsm/_0872_ heichips25_can_lehmann_fsm/_0995_ sg13g2_o21ai_1
XFILLER_21_542 VPWR VGND sg13g2_decap_8
XFILLER_21_553 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2417_ VGND VPWR heichips25_can_lehmann_fsm/_0945_ heichips25_can_lehmann_fsm/net426
+ heichips25_can_lehmann_fsm/_0108_ heichips25_can_lehmann_fsm/_0674_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2348_ heichips25_can_lehmann_fsm/net494 VPWR heichips25_can_lehmann_fsm/_0640_
+ VGND heichips25_can_lehmann_fsm/net1115 heichips25_can_lehmann_fsm/net382 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2279_ heichips25_can_lehmann_fsm/net328 VPWR heichips25_can_lehmann_fsm/_0594_
+ VGND heichips25_can_lehmann_fsm/net1191 heichips25_can_lehmann_fsm/net208 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm_fanout173 heichips25_can_lehmann_fsm/net174 heichips25_can_lehmann_fsm/net173
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout162 heichips25_can_lehmann_fsm/net163 heichips25_can_lehmann_fsm/net162
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout195 heichips25_can_lehmann_fsm/net196 heichips25_can_lehmann_fsm/net195
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout184 heichips25_can_lehmann_fsm/net187 heichips25_can_lehmann_fsm/net184
+ VPWR VGND sg13g2_buf_1
XFILLER_1_947 VPWR VGND sg13g2_decap_8
XFILLER_29_32 VPWR VGND sg13g2_decap_8
XFILLER_29_65 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2300_ heichips25_sap3/_1363_ heichips25_sap3/_1441_ heichips25_sap3/_1721_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__3280_ heichips25_sap3/_0892_ heichips25_sap3/net134 heichips25_sap3__3964_/Q
+ heichips25_sap3/net138 heichips25_sap3__3972_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2231_ heichips25_sap3/_1652_ heichips25_sap3/_1469_ heichips25_sap3/_1651_
+ VPWR VGND sg13g2_nand2_1
XFILLER_44_656 VPWR VGND sg13g2_fill_1
XFILLER_43_155 VPWR VGND sg13g2_decap_8
XFILLER_43_144 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2162_ heichips25_sap3/_1583_ heichips25_sap3/_1569_ heichips25_sap3/_1498_
+ heichips25_sap3/_1527_ heichips25_sap3/_1504_ VPWR VGND sg13g2_a22oi_1
XFILLER_31_317 VPWR VGND sg13g2_decap_8
XFILLER_32_818 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2093_ heichips25_sap3/net245 heichips25_sap3/net243 heichips25_sap3/_1514_
+ VPWR VGND sg13g2_nor2_1
XFILLER_12_520 VPWR VGND sg13g2_decap_8
XFILLER_40_884 VPWR VGND sg13g2_fill_1
XFILLER_8_524 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2995_ heichips25_sap3/_0624_ heichips25_sap3/_1760_ heichips25_sap3/_0623_
+ heichips25_sap3/_1709_ heichips25_sap3/net224 VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__1946_ VPWR heichips25_sap3/_1372_ heichips25_sap3__3966_/Q VGND
+ sg13g2_inv_1
XFILLER_20_6 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3616_ heichips25_sap3/net102 heichips25_sap3/_1061_ heichips25_sap3/_1093_
+ heichips25_sap3/_1180_ VPWR VGND sg13g2_nor3_1
Xheichips25_sap3__3547_ heichips25_sap3/_1135_ VPWR heichips25_sap3/_0096_ VGND heichips25_sap3/_1395_
+ heichips25_sap3/net56 sg13g2_o21ai_1
Xheichips25_sap3__3478_ net43 heichips25_sap3/_1076_ heichips25_sap3/_1077_ VPWR VGND
+ sg13g2_nor2_1
Xheichips25_sap3__2429_ heichips25_sap3__3895_/Q uio_out_sap3\[5\] heichips25_sap3/net215
+ heichips25_sap3/_0036_ VPWR VGND sg13g2_mux2_1
XFILLER_34_133 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__1650_ VPWR heichips25_can_lehmann_fsm/_0974_ heichips25_can_lehmann_fsm/net1198
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__1581_ VPWR heichips25_can_lehmann_fsm/_0905_ heichips25_can_lehmann_fsm/net1045
+ VGND sg13g2_inv_1
XFILLER_16_892 VPWR VGND sg13g2_decap_4
XFILLER_15_391 VPWR VGND sg13g2_decap_4
XFILLER_30_383 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2202_ heichips25_can_lehmann_fsm/net325 VPWR heichips25_can_lehmann_fsm/_0533_
+ VGND heichips25_can_lehmann_fsm/net1218 heichips25_can_lehmann_fsm/net163 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2133_ heichips25_can_lehmann_fsm/_0470_ heichips25_can_lehmann_fsm/_0471_
+ heichips25_can_lehmann_fsm/_0469_ heichips25_can_lehmann_fsm/_0472_ VPWR VGND sg13g2_nand3_1
Xheichips25_can_lehmann_fsm__2064_ VGND VPWR heichips25_can_lehmann_fsm/_1215_ heichips25_can_lehmann_fsm/_0303_
+ heichips25_can_lehmann_fsm/_0411_ heichips25_can_lehmann_fsm/_0972_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2966_ net760 VGND VPWR heichips25_can_lehmann_fsm/_0191_
+ heichips25_can_lehmann_fsm__2966_/Q clknet_leaf_19_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1917_ heichips25_can_lehmann_fsm/_1227_ heichips25_can_lehmann_fsm/_1228_
+ heichips25_can_lehmann_fsm/_1225_ heichips25_can_lehmann_fsm/_1230_ VPWR VGND heichips25_can_lehmann_fsm/_1229_
+ sg13g2_nand4_1
Xheichips25_can_lehmann_fsm__3008__530 VPWR VGND net529 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2897_ net701 VGND VPWR heichips25_can_lehmann_fsm/_0122_
+ heichips25_can_lehmann_fsm__2897_/Q clknet_leaf_21_clk sg13g2_dfrbpq_1
XFILLER_41_604 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1848_ VPWR heichips25_can_lehmann_fsm/_1164_ heichips25_can_lehmann_fsm/_1163_
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm_hold1101 heichips25_can_lehmann_fsm__2893_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1100 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__1779_ heichips25_can_lehmann_fsm/_1092_ heichips25_can_lehmann_fsm/_1093_
+ heichips25_can_lehmann_fsm/_1091_ heichips25_can_lehmann_fsm/_1095_ VPWR VGND heichips25_can_lehmann_fsm/_1094_
+ sg13g2_nand4_1
Xheichips25_can_lehmann_fsm_hold1112 heichips25_can_lehmann_fsm/_0101_ VPWR VGND heichips25_can_lehmann_fsm/net1111
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1123 heichips25_can_lehmann_fsm__3001_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1122 sg13g2_dlygate4sd3_1
XFILLER_15_78 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm_hold1134 heichips25_can_lehmann_fsm/_0284_ VPWR VGND heichips25_can_lehmann_fsm/net1133
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1156 heichips25_can_lehmann_fsm__3051_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1155 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1189 heichips25_can_lehmann_fsm__2864_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1188 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1167 heichips25_can_lehmann_fsm/_0054_ VPWR VGND heichips25_can_lehmann_fsm/net1166
+ sg13g2_dlygate4sd3_1
Xheichips25_sap3_hold832 heichips25_sap3/_0186_ VPWR VGND heichips25_sap3/net831 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1178 heichips25_can_lehmann_fsm__2886_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1177 sg13g2_dlygate4sd3_1
XFILLER_21_394 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2804__599 VPWR VGND net598 sg13g2_tiehi
Xheichips25_sap3_fanout53 heichips25_sap3/_0786_ heichips25_sap3/net53 VPWR VGND sg13g2_buf_1
Xheichips25_sap3__2780_ heichips25_sap3/_1518_ VPWR heichips25_sap3/_0425_ VGND heichips25_sap3/_1442_
+ heichips25_sap3/_1495_ sg13g2_o21ai_1
Xheichips25_sap3_fanout64 heichips25_sap3/_0444_ heichips25_sap3/net64 VPWR VGND sg13g2_buf_1
Xoutput33 net33 uio_out[6] VPWR VGND sg13g2_buf_1
Xoutput22 net22 uio_oe[3] VPWR VGND sg13g2_buf_1
Xheichips25_sap3_fanout86 heichips25_sap3/_1737_ heichips25_sap3/net86 VPWR VGND sg13g2_buf_1
X_25__511 VPWR VGND net510 sg13g2_tielo
Xheichips25_sap3_fanout75 heichips25_sap3/net76 heichips25_sap3/net75 VPWR VGND sg13g2_buf_1
Xheichips25_sap3_fanout97 heichips25_sap3/net99 heichips25_sap3/net97 VPWR VGND sg13g2_buf_1
Xheichips25_sap3__3401_ VPWR VGND heichips25_sap3__4001_/Q heichips25_sap3/net126
+ heichips25_sap3/net146 heichips25_sap3__4017_/Q heichips25_sap3/_1008_ heichips25_sap3/net116
+ sg13g2_a221oi_1
Xheichips25_sap3__3332_ heichips25_sap3/_0936_ heichips25_sap3/_0937_ heichips25_sap3/_0938_
+ heichips25_sap3/_0941_ heichips25_sap3/_0942_ VPWR VGND sg13g2_and4_1
XFILLER_17_645 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3263_ heichips25_sap3/_0876_ heichips25_sap3/net98 heichips25_sap3/_0875_
+ VPWR VGND sg13g2_nand2_1
XFILLER_44_475 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3194_ heichips25_sap3/_0803_ heichips25_sap3/_0804_ heichips25_sap3/_0805_
+ heichips25_sap3/_0806_ heichips25_sap3/_0807_ VPWR VGND sg13g2_and4_1
Xheichips25_sap3__2214_ heichips25_sap3/_1635_ heichips25_sap3/net236 heichips25_sap3/_1543_
+ VPWR VGND sg13g2_nand2b_1
Xheichips25_sap3__2145_ heichips25_sap3__4063_/Q heichips25_sap3__4064_/Q heichips25_sap3/_1566_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__2076_ heichips25_sap3/_1497_ heichips25_sap3/net246 heichips25_sap3/_1477_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__2978_ heichips25_sap3/_0613_ heichips25_sap3/net153 heichips25_sap3/_0403_
+ heichips25_sap3/net167 heichips25_sap3/net284 VPWR VGND sg13g2_a22oi_1
XFILLER_39_214 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2820_ net566 VGND VPWR heichips25_can_lehmann_fsm/net1196
+ heichips25_can_lehmann_fsm__2820_/Q clknet_leaf_8_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2751_ VGND VPWR heichips25_can_lehmann_fsm/_0857_ heichips25_can_lehmann_fsm/net425
+ heichips25_can_lehmann_fsm/_0275_ heichips25_can_lehmann_fsm/_0841_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2682_ heichips25_can_lehmann_fsm/net465 VPWR heichips25_can_lehmann_fsm/_0807_
+ VGND heichips25_can_lehmann_fsm__3016_/Q heichips25_can_lehmann_fsm/net397 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__1702_ heichips25_can_lehmann_fsm/_1026_ heichips25_can_lehmann_fsm/_1024_
+ heichips25_can_lehmann_fsm/_1025_ VPWR VGND sg13g2_nand2_1
Xheichips25_can_lehmann_fsm__1633_ VPWR heichips25_can_lehmann_fsm/_0957_ heichips25_can_lehmann_fsm/net1085
+ VGND sg13g2_inv_1
XFILLER_35_486 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1564_ VPWR heichips25_can_lehmann_fsm/_0888_ heichips25_can_lehmann_fsm/net995
+ VGND sg13g2_inv_1
XFILLER_2_519 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2116_ heichips25_can_lehmann_fsm/_0455_ heichips25_can_lehmann_fsm/net312
+ heichips25_can_lehmann_fsm__3023_/Q heichips25_can_lehmann_fsm/net313 heichips25_can_lehmann_fsm__2927_/Q
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2047_ heichips25_can_lehmann_fsm/net324 VPWR heichips25_can_lehmann_fsm/_0396_
+ VGND heichips25_can_lehmann_fsm/net1227 heichips25_can_lehmann_fsm/net177 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2988__673 VPWR VGND net672 sg13g2_tiehi
XFILLER_26_22 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2949_ net539 VGND VPWR heichips25_can_lehmann_fsm/_0174_
+ heichips25_can_lehmann_fsm__2949_/Q clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_14_604 VPWR VGND sg13g2_decap_8
XFILLER_27_987 VPWR VGND sg13g2_decap_4
XFILLER_42_957 VPWR VGND sg13g2_fill_2
XFILLER_14_615 VPWR VGND sg13g2_fill_1
XFILLER_26_88 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3950_ heichips25_sap3/net438 VGND VPWR heichips25_sap3/_0091_ heichips25_sap3__3950_/Q
+ heichips25_sap3__4014_/CLK sg13g2_dfrbpq_1
Xheichips25_sap3__2901_ heichips25_sap3/_0541_ heichips25_sap3/net154 heichips25_sap3/_0408_
+ VPWR VGND sg13g2_nand2b_1
Xheichips25_sap3__2832_ heichips25_sap3/net70 heichips25_sap3/net287 heichips25_sap3/_0475_
+ heichips25_sap3/_0041_ VPWR VGND sg13g2_a21o_1
Xheichips25_sap3__2763_ heichips25_sap3/_0409_ heichips25_sap3/_0407_ heichips25_sap3/_0408_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_can_lehmann_fsm__2856__784 VPWR VGND net783 sg13g2_tiehi
XFILLER_49_512 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2694_ heichips25_sap3/_1886_ heichips25_sap3/_1892_ heichips25_sap3/_0340_
+ VPWR VGND sg13g2_and2_1
XFILLER_49_534 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2967__757 VPWR VGND net756 sg13g2_tiehi
Xheichips25_sap3__3315_ heichips25_sap3/net48 heichips25_sap3/net52 heichips25_sap3/net59
+ heichips25_sap3/_0926_ VPWR VGND heichips25_sap3/net50 sg13g2_nand4_1
Xheichips25_sap3__3246_ heichips25_sap3/net53 heichips25_sap3/_0857_ heichips25_sap3/_0778_
+ heichips25_sap3/_0859_ VPWR VGND sg13g2_nand3_1
XFILLER_18_998 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3177_ VPWR VGND heichips25_sap3__4009_/Q heichips25_sap3/_0789_
+ heichips25_sap3/net148 heichips25_sap3__4025_/Q heichips25_sap3/_0790_ heichips25_sap3/net117
+ sg13g2_a221oi_1
Xheichips25_sap3__2128_ heichips25_sap3/net253 heichips25_sap3/_1548_ heichips25_sap3/_1549_
+ VPWR VGND sg13g2_nor2_1
XFILLER_20_629 VPWR VGND sg13g2_fill_2
XFILLER_12_180 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2059_ heichips25_sap3/_1480_ heichips25_sap3/_1463_ heichips25_sap3/_1477_
+ VPWR VGND sg13g2_nand2_1
XFILLER_8_162 VPWR VGND sg13g2_fill_2
XFILLER_8_151 VPWR VGND sg13g2_fill_2
XFILLER_8_195 VPWR VGND sg13g2_fill_2
XFILLER_8_184 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__3011__795 VPWR VGND net794 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2803_ net600 VGND VPWR heichips25_can_lehmann_fsm/_0028_
+ heichips25_can_lehmann_fsm__2803_/Q clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_36_773 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2734_ heichips25_can_lehmann_fsm/net467 VPWR heichips25_can_lehmann_fsm/_0833_
+ VGND heichips25_can_lehmann_fsm/net908 heichips25_can_lehmann_fsm/net362 sg13g2_o21ai_1
XFILLER_23_412 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2665_ VGND VPWR heichips25_can_lehmann_fsm/_0879_ heichips25_can_lehmann_fsm/net376
+ heichips25_can_lehmann_fsm/_0232_ heichips25_can_lehmann_fsm/_0798_ sg13g2_a21oi_1
XFILLER_11_607 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1616_ VPWR heichips25_can_lehmann_fsm/_0940_ heichips25_can_lehmann_fsm/net870
+ VGND sg13g2_inv_1
XFILLER_23_478 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2596_ heichips25_can_lehmann_fsm/net480 VPWR heichips25_can_lehmann_fsm/_0764_
+ VGND heichips25_can_lehmann_fsm/net972 heichips25_can_lehmann_fsm/net360 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__1547_ VPWR heichips25_can_lehmann_fsm/_0871_ heichips25_can_lehmann_fsm/net849
+ VGND sg13g2_inv_1
XFILLER_10_117 VPWR VGND sg13g2_fill_1
XFILLER_37_21 VPWR VGND sg13g2_decap_8
XFILLER_2_1021 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3100_ VGND VPWR heichips25_sap3/_0707_ heichips25_sap3/_0712_ heichips25_sap3/_0713_
+ heichips25_sap3/_0699_ sg13g2_a21oi_1
Xheichips25_sap3__3031_ heichips25_sap3/_1527_ heichips25_sap3/_1569_ heichips25_sap3/_0644_
+ VPWR VGND sg13g2_nor2_1
XFILLER_26_283 VPWR VGND sg13g2_decap_8
XFILLER_14_478 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__3023__699 VPWR VGND net698 sg13g2_tiehi
XFILLER_6_633 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3933_ heichips25_sap3/net433 VGND VPWR heichips25_sap3/_0074_ heichips25_sap3__3933_/Q
+ clkload18/A sg13g2_dfrbpq_1
XFILLER_5_143 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3864_ heichips25_sap3__3883_/Q heichips25_sap3/net1121 heichips25_sap3/net341
+ heichips25_sap3/_0191_ VPWR VGND sg13g2_mux2_1
Xheichips25_sap3__2815_ heichips25_sap3/_0458_ VPWR heichips25_sap3/_0459_ VGND heichips25_sap3/net286
+ heichips25_sap3/_0441_ sg13g2_o21ai_1
Xheichips25_sap3__3795_ heichips25_sap3/_1304_ heichips25_sap3/_1282_ heichips25_sap3__3950_/Q
+ heichips25_sap3/net292 heichips25_sap3__3958_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2746_ heichips25_sap3/_0361_ heichips25_sap3/_0391_ heichips25_sap3/_0392_
+ VPWR VGND sg13g2_nor2_1
XFILLER_49_331 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2677_ heichips25_sap3/_0329_ VPWR heichips25_sap3/_0024_ VGND heichips25_sap3/_1381_
+ heichips25_sap3/net214 sg13g2_o21ai_1
XFILLER_49_375 VPWR VGND sg13g2_decap_8
XFILLER_49_386 VPWR VGND sg13g2_fill_2
XFILLER_18_762 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3229_ heichips25_sap3/_0842_ heichips25_sap3__4004_/Q heichips25_sap3/net147
+ VPWR VGND sg13g2_nand2_1
Xheichips25_can_lehmann_fsm__2450_ heichips25_can_lehmann_fsm/net468 VPWR heichips25_can_lehmann_fsm/_0691_
+ VGND heichips25_can_lehmann_fsm/net1069 heichips25_can_lehmann_fsm/net398 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2381_ VGND VPWR heichips25_can_lehmann_fsm/_0956_ heichips25_can_lehmann_fsm/net382
+ heichips25_can_lehmann_fsm/_0090_ heichips25_can_lehmann_fsm/_0656_ sg13g2_a21oi_1
XFILLER_9_482 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm_fanout503 _00_ heichips25_can_lehmann_fsm/net503 VPWR
+ VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm__3002_ net577 VGND VPWR heichips25_can_lehmann_fsm/_0227_
+ heichips25_can_lehmann_fsm__3002_/Q clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_36_581 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2717_ VGND VPWR heichips25_can_lehmann_fsm/_0866_ heichips25_can_lehmann_fsm/net412
+ heichips25_can_lehmann_fsm/_0258_ heichips25_can_lehmann_fsm/_0824_ sg13g2_a21oi_1
XFILLER_11_415 VPWR VGND sg13g2_decap_4
XFILLER_23_253 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2648_ heichips25_can_lehmann_fsm/net472 VPWR heichips25_can_lehmann_fsm/_0790_
+ VGND heichips25_can_lehmann_fsm/net844 heichips25_can_lehmann_fsm/net404 sg13g2_o21ai_1
XFILLER_23_297 VPWR VGND sg13g2_decap_4
XFILLER_7_408 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2579_ VGND VPWR heichips25_can_lehmann_fsm/_0903_ heichips25_can_lehmann_fsm/net411
+ heichips25_can_lehmann_fsm/_0189_ heichips25_can_lehmann_fsm/_0755_ sg13g2_a21oi_1
XFILLER_3_625 VPWR VGND sg13g2_fill_2
XFILLER_3_4 VPWR VGND sg13g2_decap_8
XFILLER_2_124 VPWR VGND sg13g2_fill_1
XFILLER_2_135 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2600_ heichips25_sap3/_0272_ heichips25_sap3/_0270_ heichips25_sap3/_0271_
+ VPWR VGND sg13g2_xnor2_1
XFILLER_2_168 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2775__590 VPWR VGND net589 sg13g2_tiehi
Xheichips25_sap3__3580_ heichips25_sap3/net100 heichips25_sap3/_1157_ heichips25_sap3/_1158_
+ VPWR VGND sg13g2_nor2_1
XFILLER_48_31 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2531_ heichips25_sap3/_0208_ heichips25_sap3/net82 heichips25_sap3__3971_/Q
+ heichips25_sap3/net86 heichips25_sap3__3955_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_48_64 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2462_ heichips25_sap3/_1875_ heichips25_sap3/_1621_ heichips25_sap3/_1874_
+ VPWR VGND sg13g2_nand2_1
XFILLER_0_16 VPWR VGND sg13g2_fill_1
XFILLER_46_367 VPWR VGND sg13g2_fill_1
XFILLER_46_356 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2393_ heichips25_sap3/_1654_ heichips25_sap3/_1803_ heichips25_sap3/_1811_
+ heichips25_sap3/_1812_ VPWR VGND sg13g2_or3_1
XFILLER_34_507 VPWR VGND sg13g2_decap_8
XFILLER_15_732 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__4063_ heichips25_sap3/net433 VGND VPWR heichips25_sap3/_0003_ heichips25_sap3__4063_/Q
+ net822 sg13g2_dfrbpq_1
Xheichips25_sap3__3014_ heichips25_sap3/net233 uio_out_sap3\[2\] heichips25_sap3/_0633_
+ VPWR VGND sg13g2_nor2_1
XFILLER_9_69 VPWR VGND sg13g2_decap_8
XFILLER_11_960 VPWR VGND sg13g2_decap_4
XFILLER_6_463 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3916_ heichips25_sap3/net435 VGND VPWR heichips25_sap3/_0057_ heichips25_sap3__3916_/Q
+ heichips25_sap3__3927_/CLK sg13g2_dfrbpq_1
XFILLER_6_496 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3847_ heichips25_sap3/net838 heichips25_sap3/_1346_ heichips25_sap3/_1347_
+ VPWR VGND sg13g2_nor2_1
XFILLER_36_4 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3778_ VGND VPWR heichips25_sap3__3964_/Q heichips25_sap3/_1279_
+ heichips25_sap3/_1289_ heichips25_sap3/net290 sg13g2_a21oi_1
Xheichips25_sap3__2729_ heichips25_sap3/_0375_ heichips25_sap3/_0361_ heichips25_sap3/_0365_
+ VPWR VGND sg13g2_xnor2_1
Xheichips25_can_lehmann_fsm__1950_ heichips25_can_lehmann_fsm/_0313_ heichips25_can_lehmann_fsm/_1235_
+ heichips25_can_lehmann_fsm/_1215_ VPWR VGND sg13g2_nand2b_1
XFILLER_49_183 VPWR VGND sg13g2_decap_8
XFILLER_38_835 VPWR VGND sg13g2_fill_2
XFILLER_37_323 VPWR VGND sg13g2_decap_8
XFILLER_37_312 VPWR VGND sg13g2_fill_2
XFILLER_37_356 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1881_ heichips25_can_lehmann_fsm/net219 heichips25_can_lehmann_fsm/_1194_
+ heichips25_can_lehmann_fsm/_1195_ VPWR VGND sg13g2_nor2_1
Xheichips25_can_lehmann_fsm__2502_ heichips25_can_lehmann_fsm/net493 VPWR heichips25_can_lehmann_fsm/_0717_
+ VGND heichips25_can_lehmann_fsm__2926_/Q heichips25_can_lehmann_fsm/net405 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2433_ VGND VPWR heichips25_can_lehmann_fsm/_0939_ heichips25_can_lehmann_fsm/net370
+ heichips25_can_lehmann_fsm/_0116_ heichips25_can_lehmann_fsm/_0682_ sg13g2_a21oi_1
X_12__524 VPWR VGND net523 sg13g2_tielo
Xheichips25_can_lehmann_fsm__2364_ heichips25_can_lehmann_fsm/net500 VPWR heichips25_can_lehmann_fsm/_0648_
+ VGND heichips25_can_lehmann_fsm/net941 heichips25_can_lehmann_fsm/net387 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2295_ VGND VPWR heichips25_can_lehmann_fsm/net208 heichips25_can_lehmann_fsm/_0605_
+ heichips25_can_lehmann_fsm/_0054_ heichips25_can_lehmann_fsm/_0606_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm_fanout322 heichips25_can_lehmann_fsm/net323 heichips25_can_lehmann_fsm/net322
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout311 heichips25_can_lehmann_fsm/net312 heichips25_can_lehmann_fsm/net311
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout300 heichips25_can_lehmann_fsm/net304 heichips25_can_lehmann_fsm/net300
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout344 heichips25_can_lehmann_fsm__2800_/Q heichips25_can_lehmann_fsm/net344
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout333 heichips25_can_lehmann_fsm/net334 heichips25_can_lehmann_fsm/net333
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout355 heichips25_can_lehmann_fsm/net356 heichips25_can_lehmann_fsm/net355
+ VPWR VGND sg13g2_buf_1
Xclkbuf_5_4__f_heichips25_sap3\_sap_3_inst.alu_inst.clk heichips25_sap3__4012_/CLK
+ clknet_4_2_0_heichips25_sap3\/sap_3_inst.alu_inst.clk VPWR VGND sg13g2_buf_16
Xheichips25_can_lehmann_fsm_fanout366 heichips25_can_lehmann_fsm/net367 heichips25_can_lehmann_fsm/net366
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout388 heichips25_can_lehmann_fsm/net389 heichips25_can_lehmann_fsm/net388
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout399 heichips25_can_lehmann_fsm/net400 heichips25_can_lehmann_fsm/net399
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout377 heichips25_can_lehmann_fsm/net379 heichips25_can_lehmann_fsm/net377
+ VPWR VGND sg13g2_buf_1
XFILLER_28_334 VPWR VGND sg13g2_fill_1
XFILLER_43_315 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__1962_ VPWR heichips25_sap3/_1388_ heichips25_sap3__3980_/Q VGND
+ sg13g2_inv_1
Xheichips25_sap3__3701_ heichips25_sap3/_1231_ VPWR heichips25_sap3/_0152_ VGND heichips25_sap3/_1232_
+ heichips25_sap3/_1233_ sg13g2_o21ai_1
Xheichips25_sap3__3632_ heichips25_sap3/_1189_ heichips25_sap3/_1188_ heichips25_sap3/_1056_
+ heichips25_sap3/net93 heichips25_sap3__3987_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_3_499 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3563_ heichips25_sap3/_1144_ heichips25_sap3/net134 heichips25_sap3/net131
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__2514_ heichips25_sap3__3892_/Q VPWR heichips25_sap3/_1925_ VGND
+ heichips25_sap3/_1717_ heichips25_sap3/_1878_ sg13g2_o21ai_1
XFILLER_47_621 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2814__579 VPWR VGND net578 sg13g2_tiehi
Xheichips25_sap3__3494_ heichips25_sap3/net108 heichips25_sap3/_1054_ heichips25_sap3/_1091_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__2445_ VPWR VGND heichips25_sap3__3983_/Q heichips25_sap3/net80 heichips25_sap3/net72
+ heichips25_sap3__4015_/Q heichips25_sap3/_1860_ heichips25_sap3/net217 sg13g2_a221oi_1
XFILLER_19_356 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2376_ heichips25_sap3/_1797_ heichips25_sap3/net73 heichips25_sap3__4010_/Q
+ heichips25_sap3/net90 heichips25_sap3__3946_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_35_816 VPWR VGND sg13g2_decap_8
XFILLER_34_315 VPWR VGND sg13g2_decap_4
XFILLER_34_359 VPWR VGND sg13g2_fill_1
XFILLER_15_562 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__4046_ heichips25_sap3/net452 VGND VPWR heichips25_sap3/_0187_ heichips25_sap3__4046_/Q
+ clknet_leaf_22_clk sg13g2_dfrbpq_1
XFILLER_7_761 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2080_ VPWR VGND heichips25_can_lehmann_fsm/_0423_ heichips25_can_lehmann_fsm/net182
+ heichips25_can_lehmann_fsm/net186 heichips25_can_lehmann_fsm/net345 heichips25_can_lehmann_fsm/_0424_
+ heichips25_can_lehmann_fsm/net190 sg13g2_a221oi_1
XFILLER_38_610 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2982_ net696 VGND VPWR heichips25_can_lehmann_fsm/_0207_
+ heichips25_can_lehmann_fsm__2982_/Q clknet_leaf_14_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1933_ heichips25_can_lehmann_fsm/net337 VPWR heichips25_can_lehmann_fsm/_0296_
+ VGND heichips25_can_lehmann_fsm__2978_/Q heichips25_can_lehmann_fsm/net338 sg13g2_o21ai_1
XFILLER_38_698 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1864_ heichips25_can_lehmann_fsm/_1179_ heichips25_can_lehmann_fsm/net332
+ heichips25_can_lehmann_fsm__3035_/Q heichips25_can_lehmann_fsm/net307 heichips25_can_lehmann_fsm__2939_/Q
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3_fanout204 heichips25_sap3/_0436_ heichips25_sap3/net204 VPWR VGND
+ sg13g2_buf_1
X_29_ net514 uio_oe_sap3\[7\] net506 net26 VPWR VGND sg13g2_mux2_1
Xheichips25_sap3_fanout248 heichips25_sap3/_1453_ heichips25_sap3/net248 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout226 heichips25_sap3/_1598_ heichips25_sap3/net226 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout215 heichips25_sap3/_1801_ heichips25_sap3/net215 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout237 heichips25_sap3/net239 heichips25_sap3/net237 VPWR VGND
+ sg13g2_buf_1
XFILLER_40_307 VPWR VGND sg13g2_fill_2
Xheichips25_sap3_fanout259 heichips25_sap3__3930_/Q heichips25_sap3/net259 VPWR VGND
+ sg13g2_buf_1
Xheichips25_can_lehmann_fsm__1795_ VPWR VGND heichips25_can_lehmann_fsm__2973_/Q heichips25_can_lehmann_fsm/_1110_
+ heichips25_can_lehmann_fsm/net294 heichips25_can_lehmann_fsm__2949_/Q heichips25_can_lehmann_fsm/_1111_
+ heichips25_can_lehmann_fsm/net306 sg13g2_a221oi_1
Xheichips25_can_lehmann_fsm__2416_ heichips25_can_lehmann_fsm/net499 VPWR heichips25_can_lehmann_fsm/_0674_
+ VGND heichips25_can_lehmann_fsm__2883_/Q heichips25_can_lehmann_fsm/net426 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2347_ VGND VPWR heichips25_can_lehmann_fsm/_0965_ heichips25_can_lehmann_fsm/net406
+ heichips25_can_lehmann_fsm/_0073_ heichips25_can_lehmann_fsm/_0639_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2278_ VGND VPWR heichips25_can_lehmann_fsm/net968 heichips25_can_lehmann_fsm/net172
+ heichips25_can_lehmann_fsm/_0593_ heichips25_can_lehmann_fsm/_0592_ sg13g2_a21oi_1
XFILLER_20_35 VPWR VGND sg13g2_fill_2
XFILLER_20_68 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm_fanout174 heichips25_can_lehmann_fsm/_0557_ heichips25_can_lehmann_fsm/net174
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout163 heichips25_can_lehmann_fsm/_0498_ heichips25_can_lehmann_fsm/net163
+ VPWR VGND sg13g2_buf_1
XFILLER_1_926 VPWR VGND sg13g2_decap_8
XFILLER_49_908 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_fanout196 heichips25_can_lehmann_fsm/_0306_ heichips25_can_lehmann_fsm/net196
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout185 heichips25_can_lehmann_fsm/net187 heichips25_can_lehmann_fsm/net185
+ VPWR VGND sg13g2_buf_1
XFILLER_29_88 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2230_ heichips25_sap3/net227 heichips25_sap3/_1613_ heichips25_sap3/_1651_
+ VPWR VGND sg13g2_and2_1
XFILLER_16_304 VPWR VGND sg13g2_fill_1
XFILLER_28_164 VPWR VGND sg13g2_decap_4
XFILLER_43_134 VPWR VGND sg13g2_decap_4
XFILLER_43_101 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2161_ heichips25_sap3/net245 VPWR heichips25_sap3/_1582_ VGND heichips25_sap3/_1499_
+ heichips25_sap3/_1581_ sg13g2_o21ai_1
XFILLER_25_860 VPWR VGND sg13g2_decap_4
XFILLER_43_178 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2092_ heichips25_sap3/net257 heichips25_sap3/_1438_ heichips25_sap3/net255
+ heichips25_sap3/_1511_ heichips25_sap3/_1513_ VPWR VGND sg13g2_or4_1
XFILLER_24_370 VPWR VGND sg13g2_fill_2
Xclkbuf_4_1_0_heichips25_sap3\_sap_3_inst.alu_inst.clk clknet_0_heichips25_sap3\/sap_3_inst.alu_inst.clk
+ clknet_4_1_0_heichips25_sap3\/sap_3_inst.alu_inst.clk VPWR VGND sg13g2_buf_8
XFILLER_6_48 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2994_ VGND VPWR heichips25_sap3/net238 heichips25_sap3/_1614_ heichips25_sap3/_0623_
+ heichips25_sap3/_1662_ sg13g2_a21oi_1
XFILLER_6_59 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__1945_ VPWR heichips25_sap3/_1371_ heichips25_sap3__3982_/Q VGND
+ sg13g2_inv_1
Xheichips25_sap3__3615_ heichips25_sap3/_1179_ VPWR heichips25_sap3/_0120_ VGND heichips25_sap3/_1394_
+ heichips25_sap3/net141 sg13g2_o21ai_1
XFILLER_0_992 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3546_ heichips25_sap3/_1057_ heichips25_sap3/net56 heichips25_sap3/_1056_
+ heichips25_sap3/_1135_ VPWR VGND sg13g2_nand3_1
Xheichips25_sap3__3477_ heichips25_sap3/net121 heichips25_sap3/_1025_ heichips25_sap3/_1076_
+ VPWR VGND sg13g2_and2_1
Xheichips25_sap3__2428_ heichips25_sap3/_1831_ heichips25_sap3/_1836_ heichips25_sap3/_1844_
+ uio_out_sap3\[5\] VPWR VGND sg13g2_or3_1
Xheichips25_can_lehmann_fsm__2866__764 VPWR VGND net763 sg13g2_tiehi
Xheichips25_sap3__2359_ heichips25_sap3/_1780_ heichips25_sap3/_1775_ heichips25_sap3/_1779_
+ VPWR VGND sg13g2_nand2_1
XFILLER_16_860 VPWR VGND sg13g2_fill_1
XFILLER_34_145 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1580_ VPWR heichips25_can_lehmann_fsm/_0904_ heichips25_can_lehmann_fsm/net1017
+ VGND sg13g2_inv_1
XFILLER_22_318 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__4029_ heichips25_sap3/net461 VGND VPWR heichips25_sap3/_0170_ heichips25_sap3__4029_/Q
+ clknet_leaf_2_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2201_ heichips25_can_lehmann_fsm/_0532_ heichips25_can_lehmann_fsm/net165
+ heichips25_can_lehmann_fsm/_0531_ heichips25_can_lehmann_fsm/net175 heichips25_can_lehmann_fsm/net974
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2132_ heichips25_can_lehmann_fsm/_0471_ heichips25_can_lehmann_fsm/net307
+ heichips25_can_lehmann_fsm__2958_/Q heichips25_can_lehmann_fsm/net315 heichips25_can_lehmann_fsm__2934_/Q
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2063_ VPWR VGND heichips25_can_lehmann_fsm/net195 heichips25_can_lehmann_fsm/_0410_
+ heichips25_can_lehmann_fsm/_0408_ heichips25_can_lehmann_fsm/_0398_ heichips25_can_lehmann_fsm/_0018_
+ heichips25_can_lehmann_fsm/_0407_ sg13g2_a221oi_1
Xheichips25_can_lehmann_fsm__3014__771 VPWR VGND net770 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2965_ net764 VGND VPWR heichips25_can_lehmann_fsm/net875
+ heichips25_can_lehmann_fsm__2965_/Q clknet_leaf_18_clk sg13g2_dfrbpq_1
XFILLER_39_985 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1916_ heichips25_can_lehmann_fsm/_1229_ heichips25_can_lehmann_fsm/net311
+ heichips25_can_lehmann_fsm__3027_/Q heichips25_can_lehmann_fsm/net318 heichips25_can_lehmann_fsm__3003_/Q
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2896_ net703 VGND VPWR heichips25_can_lehmann_fsm/_0121_
+ heichips25_can_lehmann_fsm__2896_/Q clknet_leaf_22_clk sg13g2_dfrbpq_1
XFILLER_25_101 VPWR VGND sg13g2_decap_4
XFILLER_26_657 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1847_ heichips25_can_lehmann_fsm/_1139_ heichips25_can_lehmann_fsm/_1161_
+ heichips25_can_lehmann_fsm/_1163_ VPWR VGND sg13g2_nor2_1
XFILLER_41_638 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1778_ VGND VPWR heichips25_can_lehmann_fsm__3013_/Q heichips25_can_lehmann_fsm/net310
+ heichips25_can_lehmann_fsm/_1094_ heichips25_can_lehmann_fsm/net302 sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm_hold1102 heichips25_can_lehmann_fsm/_0119_ VPWR VGND heichips25_can_lehmann_fsm/net1101
+ sg13g2_dlygate4sd3_1
XFILLER_13_318 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm_hold1124 heichips25_can_lehmann_fsm/_0226_ VPWR VGND heichips25_can_lehmann_fsm/net1123
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1157 heichips25_can_lehmann_fsm/_0277_ VPWR VGND heichips25_can_lehmann_fsm/net1156
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1135 heichips25_can_lehmann_fsm__3002_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1134 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__2960__785 VPWR VGND net784 sg13g2_tiehi
Xheichips25_can_lehmann_fsm_hold1168 heichips25_can_lehmann_fsm__2871_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1167 sg13g2_dlygate4sd3_1
Xheichips25_sap3_hold833 heichips25_sap3__4062_/Q VPWR VGND heichips25_sap3/net832
+ sg13g2_dlygate4sd3_1
XFILLER_31_34 VPWR VGND sg13g2_decap_8
Xheichips25_sap3_fanout54 heichips25_sap3/_0786_ heichips25_sap3/net54 VPWR VGND sg13g2_buf_1
Xheichips25_sap3_fanout87 heichips25_sap3/net88 heichips25_sap3/net87 VPWR VGND sg13g2_buf_1
Xheichips25_sap3_fanout65 heichips25_sap3/_0444_ heichips25_sap3/net65 VPWR VGND sg13g2_buf_1
Xoutput34 net34 uio_out[7] VPWR VGND sg13g2_buf_1
Xoutput23 net23 uio_oe[4] VPWR VGND sg13g2_buf_1
Xheichips25_sap3_fanout76 heichips25_sap3/_1744_ heichips25_sap3/net76 VPWR VGND sg13g2_buf_1
Xheichips25_sap3_fanout98 heichips25_sap3/net99 heichips25_sap3/net98 VPWR VGND sg13g2_buf_1
XFILLER_49_716 VPWR VGND sg13g2_decap_8
XFILLER_49_738 VPWR VGND sg13g2_fill_2
XFILLER_49_727 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3400_ heichips25_sap3/_0077_ heichips25_sap3/_0997_ heichips25_sap3/_1007_
+ heichips25_sap3/net55 heichips25_sap3/_1404_ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3331_ heichips25_sap3/_0939_ heichips25_sap3/_0940_ heichips25_sap3/_0941_
+ VPWR VGND sg13g2_and2_1
Xheichips25_sap3__3262_ heichips25_sap3/net49 heichips25_sap3/net59 heichips25_sap3/_0874_
+ heichips25_sap3/_0875_ VPWR VGND sg13g2_a21o_1
Xheichips25_sap3__3193_ heichips25_sap3/_0717_ heichips25_sap3/net151 heichips25_sap3__4023_/Q
+ heichips25_sap3/_0806_ VPWR VGND sg13g2_nand3_1
Xheichips25_sap3__2213_ heichips25_sap3/_1630_ heichips25_sap3/_1631_ heichips25_sap3/_1612_
+ heichips25_sap3/_1634_ VPWR VGND heichips25_sap3/_1633_ sg13g2_nand4_1
XFILLER_17_668 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__3026__675 VPWR VGND net674 sg13g2_tiehi
Xheichips25_sap3__2144_ heichips25_sap3/net257 heichips25_sap3/net269 heichips25_sap3/_1565_
+ VPWR VGND heichips25_sap3/_1529_ sg13g2_nand3b_1
Xclkbuf_5_22__f_heichips25_sap3\_sap_3_inst.alu_inst.clk heichips25_sap3__3920_/CLK
+ clknet_4_11_0_heichips25_sap3\/sap_3_inst.alu_inst.clk VPWR VGND sg13g2_buf_16
XFILLER_25_690 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2075_ heichips25_sap3/net246 heichips25_sap3/_1477_ heichips25_sap3/_1496_
+ VPWR VGND sg13g2_and2_1
XFILLER_8_344 VPWR VGND sg13g2_decap_8
XFILLER_9_878 VPWR VGND sg13g2_fill_2
XFILLER_12_373 VPWR VGND sg13g2_fill_2
XFILLER_12_395 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2977_ heichips25_sap3/_0612_ heichips25_sap3__3909_/Q heichips25_sap3/_0607_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__3529_ heichips25_sap3/_1121_ heichips25_sap3/net97 heichips25_sap3/_0994_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_can_lehmann_fsm__2750_ heichips25_can_lehmann_fsm/net491 VPWR heichips25_can_lehmann_fsm/_0841_
+ VGND heichips25_can_lehmann_fsm__3050_/Q heichips25_can_lehmann_fsm/net425 sg13g2_o21ai_1
XFILLER_36_933 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1701_ VGND VPWR heichips25_can_lehmann_fsm__3039_/Q heichips25_can_lehmann_fsm/net331
+ heichips25_can_lehmann_fsm/_1025_ heichips25_can_lehmann_fsm/net300 sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2681_ VGND VPWR heichips25_can_lehmann_fsm/_0875_ heichips25_can_lehmann_fsm/net358
+ heichips25_can_lehmann_fsm/_0240_ heichips25_can_lehmann_fsm/_0806_ sg13g2_a21oi_1
XFILLER_23_605 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1632_ VPWR heichips25_can_lehmann_fsm/_0956_ heichips25_can_lehmann_fsm/net883
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__1563_ VPWR heichips25_can_lehmann_fsm/_0887_ heichips25_can_lehmann_fsm/net928
+ VGND sg13g2_inv_1
XFILLER_22_126 VPWR VGND sg13g2_decap_8
XFILLER_31_671 VPWR VGND sg13g2_fill_1
XFILLER_7_91 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2115_ heichips25_can_lehmann_fsm/_0454_ heichips25_can_lehmann_fsm/net331
+ heichips25_can_lehmann_fsm__3047_/Q heichips25_can_lehmann_fsm/net306 heichips25_can_lehmann_fsm__2951_/Q
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2046_ heichips25_can_lehmann_fsm/_0394_ heichips25_can_lehmann_fsm/_0391_
+ heichips25_can_lehmann_fsm/_0393_ heichips25_can_lehmann_fsm/_0395_ VPWR VGND sg13g2_a21o_1
XFILLER_45_207 VPWR VGND sg13g2_decap_8
XFILLER_38_281 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2948_ net543 VGND VPWR heichips25_can_lehmann_fsm/_0173_
+ heichips25_can_lehmann_fsm__2948_/Q clknet_leaf_0_clk sg13g2_dfrbpq_1
XFILLER_42_903 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2879_ net737 VGND VPWR heichips25_can_lehmann_fsm/_0104_
+ heichips25_can_lehmann_fsm__2879_/Q clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_42_947 VPWR VGND sg13g2_fill_1
XFILLER_41_413 VPWR VGND sg13g2_fill_2
XFILLER_14_649 VPWR VGND sg13g2_fill_1
XFILLER_6_826 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2900_ heichips25_sap3/_0540_ heichips25_sap3/_0449_ heichips25_sap3/_0351_
+ heichips25_sap3/_0445_ heichips25_sap3/_0380_ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2995__634 VPWR VGND net633 sg13g2_tiehi
XFILLER_5_325 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2831_ VPWR VGND heichips25_sap3/_0474_ heichips25_sap3/net70 heichips25_sap3/_0473_
+ heichips25_sap3/_1922_ heichips25_sap3/_0475_ heichips25_sap3/net158 sg13g2_a221oi_1
Xheichips25_sap3__2762_ heichips25_sap3/_0408_ heichips25_sap3/_0380_ heichips25_sap3/_0396_
+ VPWR VGND sg13g2_xnor2_1
Xheichips25_sap3__2693_ VGND VPWR heichips25_sap3/_0339_ heichips25_sap3/_0337_ heichips25_sap3/_1887_
+ sg13g2_or2_1
Xheichips25_sap3__3314_ heichips25_sap3/_0924_ VPWR heichips25_sap3/_0925_ VGND heichips25_sap3/net127
+ heichips25_sap3/_0914_ sg13g2_o21ai_1
XFILLER_18_966 VPWR VGND sg13g2_fill_2
XFILLER_18_977 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3245_ heichips25_sap3/net53 heichips25_sap3/_0857_ heichips25_sap3/_0858_
+ VPWR VGND sg13g2_and2_1
Xheichips25_sap3__3176_ heichips25_sap3/_0789_ heichips25_sap3/_0787_ heichips25_sap3/_0788_
+ VPWR VGND sg13g2_nand2_1
XFILLER_41_980 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2127_ heichips25_sap3__4066_/Q heichips25_sap3/net252 heichips25_sap3/_1548_
+ VPWR VGND heichips25_sap3__4065_/Q sg13g2_nand3b_1
Xheichips25_sap3__2058_ heichips25_sap3/_1464_ heichips25_sap3/_1478_ heichips25_sap3/_1479_
+ VPWR VGND sg13g2_nor2_1
XFILLER_12_192 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2974__729 VPWR VGND net728 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2802_ net602 VGND VPWR heichips25_can_lehmann_fsm/_0027_
+ heichips25_can_lehmann_fsm__2802_/Q clknet_leaf_5_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2733_ VGND VPWR heichips25_can_lehmann_fsm/_0862_ heichips25_can_lehmann_fsm/net393
+ heichips25_can_lehmann_fsm/_0266_ heichips25_can_lehmann_fsm/_0832_ sg13g2_a21oi_1
XFILLER_35_251 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2664_ heichips25_can_lehmann_fsm/net487 VPWR heichips25_can_lehmann_fsm/_0798_
+ VGND heichips25_can_lehmann_fsm__3006_/Q heichips25_can_lehmann_fsm/net376 sg13g2_o21ai_1
XFILLER_35_295 VPWR VGND sg13g2_decap_8
XFILLER_23_446 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1615_ VPWR heichips25_can_lehmann_fsm/_0939_ heichips25_can_lehmann_fsm/net955
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__2595_ VGND VPWR heichips25_can_lehmann_fsm/_0899_ heichips25_can_lehmann_fsm/net400
+ heichips25_can_lehmann_fsm/_0197_ heichips25_can_lehmann_fsm/_0763_ sg13g2_a21oi_1
XFILLER_23_468 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1546_ VPWR heichips25_can_lehmann_fsm/_0870_ heichips25_can_lehmann_fsm/net1074
+ VGND sg13g2_inv_1
XFILLER_12_69 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2029_ heichips25_can_lehmann_fsm/_0380_ heichips25_can_lehmann_fsm/_0980_
+ heichips25_can_lehmann_fsm/_1071_ VPWR VGND sg13g2_xnor2_1
XFILLER_37_55 VPWR VGND sg13g2_decap_4
XFILLER_37_44 VPWR VGND sg13g2_decap_4
XFILLER_2_1000 VPWR VGND sg13g2_decap_8
XFILLER_18_218 VPWR VGND sg13g2_decap_8
XFILLER_27_763 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3030_ VGND VPWR heichips25_sap3/_1485_ heichips25_sap3/_0642_ heichips25_sap3/_0643_
+ heichips25_sap3/_1697_ sg13g2_a21oi_1
XFILLER_41_243 VPWR VGND sg13g2_fill_1
XFILLER_14_457 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_21_clk clknet_2_0__leaf_clk clknet_leaf_21_clk VPWR VGND sg13g2_buf_8
Xheichips25_sap3__3932_ heichips25_sap3/net434 VGND VPWR heichips25_sap3/_0073_ heichips25_sap3__3932_/Q
+ heichips25_sap3__4012_/CLK sg13g2_dfrbpq_1
XFILLER_10_685 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3863_ heichips25_sap3__3882_/Q heichips25_sap3/net1145 heichips25_sap3/net341
+ heichips25_sap3/_0190_ VPWR VGND sg13g2_mux2_1
Xheichips25_sap3__2814_ heichips25_sap3/net159 VPWR heichips25_sap3/_0458_ VGND heichips25_sap3/net286
+ heichips25_sap3__3916_/Q sg13g2_o21ai_1
Xheichips25_sap3__3794_ heichips25_sap3/_1303_ heichips25_sap3/_1281_ heichips25_sap3__4014_/Q
+ heichips25_sap3/_1270_ heichips25_sap3__4022_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2745_ VGND VPWR heichips25_sap3/net286 heichips25_sap3/_1396_ heichips25_sap3/_0391_
+ heichips25_sap3/_0390_ sg13g2_a21oi_1
XFILLER_2_884 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2676_ heichips25_sap3/_0329_ heichips25_sap3__3883_/Q heichips25_sap3/net214
+ VPWR VGND sg13g2_nand2_1
XFILLER_49_354 VPWR VGND sg13g2_decap_8
XFILLER_18_785 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3228_ heichips25_sap3/_0835_ heichips25_sap3/_0840_ heichips25_sap3/_0841_
+ VPWR VGND sg13g2_and2_1
XFILLER_33_744 VPWR VGND sg13g2_decap_8
XFILLER_33_755 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3159_ heichips25_sap3/_0696_ heichips25_sap3/_0759_ heichips25_sap3/_0772_
+ VPWR VGND sg13g2_and2_1
Xheichips25_can_lehmann_fsm__2824__559 VPWR VGND net558 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2380_ heichips25_can_lehmann_fsm/net495 VPWR heichips25_can_lehmann_fsm/_0656_
+ VGND heichips25_can_lehmann_fsm__2864_/Q heichips25_can_lehmann_fsm/net382 sg13g2_o21ai_1
XFILLER_32_276 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_12_clk clknet_2_3__leaf_clk clknet_leaf_12_clk VPWR VGND sg13g2_buf_8
Xheichips25_can_lehmann_fsm__3001_ net585 VGND VPWR heichips25_can_lehmann_fsm/net1123
+ heichips25_can_lehmann_fsm__3001_/Q clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_4_92 VPWR VGND sg13g2_decap_8
XFILLER_36_560 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2716_ heichips25_can_lehmann_fsm/net484 VPWR heichips25_can_lehmann_fsm/_0824_
+ VGND heichips25_can_lehmann_fsm__3033_/Q heichips25_can_lehmann_fsm/net411 sg13g2_o21ai_1
XFILLER_24_755 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2647_ VGND VPWR heichips25_can_lehmann_fsm/_0885_ heichips25_can_lehmann_fsm/net404
+ heichips25_can_lehmann_fsm/_0223_ heichips25_can_lehmann_fsm/_0789_ sg13g2_a21oi_1
XFILLER_23_35 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2578_ heichips25_can_lehmann_fsm/net478 VPWR heichips25_can_lehmann_fsm/_0755_
+ VGND heichips25_can_lehmann_fsm/net1091 heichips25_can_lehmann_fsm/net411 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__1529_ VPWR heichips25_can_lehmann_fsm/_0853_ heichips25_can_lehmann_fsm/net1142
+ VGND sg13g2_inv_1
XFILLER_2_158 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3876__821 VPWR net820 clkload27/A VGND sg13g2_inv_1
Xheichips25_sap3__2530_ heichips25_sap3/_0207_ heichips25_sap3/net76 heichips25_sap3__3987_/Q
+ heichips25_sap3/net83 heichips25_sap3__3963_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2461_ heichips25_sap3/_1874_ heichips25_sap3/_1782_ heichips25_sap3/_1361_
+ heichips25_sap3/_1614_ heichips25_sap3/net228 VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2392_ heichips25_sap3/_1808_ heichips25_sap3/_1810_ heichips25_sap3/_1811_
+ VPWR VGND sg13g2_nor2_1
XFILLER_15_722 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__4062_ heichips25_sap3/net458 VGND VPWR heichips25_sap3__4062_/D
+ heichips25_sap3__4062_/Q clknet_leaf_1_clk sg13g2_dfrbpq_1
XFILLER_9_15 VPWR VGND sg13g2_fill_2
XFILLER_9_26 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3013_ heichips25_sap3/_0632_ VPWR heichips25_sap3/_0065_ VGND heichips25_sap3/net233
+ heichips25_sap3/_1922_ sg13g2_o21ai_1
XFILLER_30_703 VPWR VGND sg13g2_fill_2
XFILLER_14_287 VPWR VGND sg13g2_decap_8
XFILLER_14_298 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3915_ heichips25_sap3/net450 VGND VPWR heichips25_sap3/_0056_ heichips25_sap3__3915_/Q
+ heichips25_sap3__3922_/CLK sg13g2_dfrbpq_1
Xheichips25_sap3__3846_ heichips25_sap3/_0288_ VPWR heichips25_sap3/_1346_ VGND heichips25_sap3/net1225
+ heichips25_sap3/_1366_ sg13g2_o21ai_1
Xheichips25_sap3__3777_ heichips25_sap3/_1288_ heichips25_sap3/_1282_ heichips25_sap3__3948_/Q
+ heichips25_sap3/_1265_ heichips25_sap3__3996_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2728_ heichips25_sap3/_0363_ heichips25_sap3/_0372_ heichips25_sap3/net254
+ heichips25_sap3/_0374_ VPWR VGND sg13g2_nand3_1
Xheichips25_sap3__2659_ heichips25_sap3/_1468_ heichips25_sap3/_0324_ heichips25_sap3/_0004_
+ VPWR VGND sg13g2_and2_1
XFILLER_29_4 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_1_clk clknet_2_0__leaf_clk clknet_leaf_1_clk VPWR VGND sg13g2_buf_8
XFILLER_49_151 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1880_ heichips25_can_lehmann_fsm/_1193_ VPWR heichips25_can_lehmann_fsm/_1194_
+ VGND heichips25_can_lehmann_fsm/net1272 heichips25_can_lehmann_fsm/net335 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2501_ VGND VPWR heichips25_can_lehmann_fsm/_0922_ heichips25_can_lehmann_fsm/net359
+ heichips25_can_lehmann_fsm/_0150_ heichips25_can_lehmann_fsm/_0716_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2432_ heichips25_can_lehmann_fsm/net477 VPWR heichips25_can_lehmann_fsm/_0682_
+ VGND heichips25_can_lehmann_fsm__2890_/Q heichips25_can_lehmann_fsm/net370 sg13g2_o21ai_1
XFILLER_20_257 VPWR VGND sg13g2_decap_8
XFILLER_21_769 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2363_ VGND VPWR heichips25_can_lehmann_fsm/_0961_ heichips25_can_lehmann_fsm/net430
+ heichips25_can_lehmann_fsm/_0081_ heichips25_can_lehmann_fsm/_0647_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2294_ heichips25_can_lehmann_fsm/net328 VPWR heichips25_can_lehmann_fsm/_0606_
+ VGND heichips25_can_lehmann_fsm/net1165 heichips25_can_lehmann_fsm/net208 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm_fanout323 heichips25_can_lehmann_fsm/net324 heichips25_can_lehmann_fsm/net323
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout312 heichips25_can_lehmann_fsm/_0994_ heichips25_can_lehmann_fsm/net312
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout301 heichips25_can_lehmann_fsm/net304 heichips25_can_lehmann_fsm/net301
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm__2876__744 VPWR VGND net743 sg13g2_tiehi
Xheichips25_can_lehmann_fsm_fanout345 heichips25_can_lehmann_fsm/net1264 heichips25_can_lehmann_fsm/net345
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout356 heichips25_can_lehmann_fsm/net362 heichips25_can_lehmann_fsm/net356
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout334 heichips25_can_lehmann_fsm/_1003_ heichips25_can_lehmann_fsm/net334
+ VPWR VGND sg13g2_buf_1
XFILLER_47_1023 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm_fanout389 heichips25_can_lehmann_fsm/_0624_ heichips25_can_lehmann_fsm/net389
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout378 heichips25_can_lehmann_fsm/net379 heichips25_can_lehmann_fsm/net378
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout367 heichips25_can_lehmann_fsm/net389 heichips25_can_lehmann_fsm/net367
+ VPWR VGND sg13g2_buf_1
XFILLER_28_302 VPWR VGND sg13g2_decap_8
XFILLER_29_858 VPWR VGND sg13g2_fill_1
XFILLER_11_224 VPWR VGND sg13g2_fill_1
XFILLER_11_279 VPWR VGND sg13g2_fill_2
Xclkload0 clknet_leaf_0_clk clkload0/Y VPWR VGND sg13g2_inv_4
Xheichips25_sap3__1961_ VPWR heichips25_sap3/_1387_ heichips25_sap3__3996_/Q VGND
+ sg13g2_inv_1
Xheichips25_sap3__3700_ uio_oe_sap3\[0\] heichips25_sap3/_1055_ heichips25_sap3/_1086_
+ heichips25_sap3/_1233_ VPWR VGND sg13g2_nor3_1
XFILLER_3_434 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2777__653 VPWR VGND net652 sg13g2_tiehi
XFILLER_3_478 VPWR VGND sg13g2_decap_8
XFILLER_3_456 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3631_ VGND VPWR heichips25_sap3/net60 heichips25_sap3/net99 heichips25_sap3/_1188_
+ heichips25_sap3/net93 sg13g2_a21oi_1
Xheichips25_sap3__3562_ heichips25_sap3/_1143_ heichips25_sap3/net134 heichips25_sap3/_0876_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__2513_ heichips25_sap3/_1900_ VPWR heichips25_sap3/_0034_ VGND heichips25_sap3/_1923_
+ heichips25_sap3/_1924_ sg13g2_o21ai_1
Xheichips25_sap3__3493_ VGND VPWR heichips25_sap3/_0212_ heichips25_sap3/_1088_ heichips25_sap3/_1090_
+ heichips25_sap3/_1089_ sg13g2_a21oi_1
Xheichips25_sap3__2444_ heichips25_sap3/_1857_ heichips25_sap3/_1858_ heichips25_sap3/_1859_
+ VPWR VGND sg13g2_and2_1
Xheichips25_sap3__2375_ VPWR VGND heichips25_sap3__3970_/Q heichips25_sap3/net79 heichips25_sap3/net84
+ heichips25_sap3__4018_/Q heichips25_sap3/_1796_ heichips25_sap3/net216 sg13g2_a221oi_1
XFILLER_46_198 VPWR VGND sg13g2_fill_1
XFILLER_46_187 VPWR VGND sg13g2_fill_1
XFILLER_34_338 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__4045_ heichips25_sap3/net453 VGND VPWR heichips25_sap3/net831 heichips25_sap3__4072_/A
+ clknet_leaf_22_clk sg13g2_dfrbpq_1
XFILLER_42_382 VPWR VGND sg13g2_fill_1
XFILLER_15_585 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_hold990 heichips25_can_lehmann_fsm__2892_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net989 sg13g2_dlygate4sd3_1
XFILLER_7_795 VPWR VGND sg13g2_decap_8
XFILLER_7_784 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3829_ heichips25_sap3/net340 heichips25_sap3/net953 heichips25_sap3/_1334_
+ heichips25_sap3/_0179_ VPWR VGND sg13g2_a21o_1
Xheichips25_can_lehmann_fsm__2981_ net700 VGND VPWR heichips25_can_lehmann_fsm/net1023
+ heichips25_can_lehmann_fsm__2981_/Q clknet_leaf_14_clk sg13g2_dfrbpq_1
XFILLER_37_121 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__1932_ heichips25_can_lehmann_fsm/_0295_ heichips25_can_lehmann_fsm__2906_/Q
+ heichips25_can_lehmann_fsm/net298 VPWR VGND sg13g2_nand2_1
XFILLER_38_688 VPWR VGND sg13g2_fill_1
X_28_ net513 uio_oe_sap3\[6\] net506 net25 VPWR VGND sg13g2_mux2_1
Xheichips25_can_lehmann_fsm__1863_ VGND VPWR heichips25_can_lehmann_fsm__2987_/Q heichips25_can_lehmann_fsm/net318
+ heichips25_can_lehmann_fsm/_1178_ heichips25_can_lehmann_fsm/net302 sg13g2_a21oi_1
Xheichips25_sap3_fanout227 heichips25_sap3/net228 heichips25_sap3/net227 VPWR VGND
+ sg13g2_buf_1
XFILLER_1_93 VPWR VGND sg13g2_decap_4
Xheichips25_sap3_fanout238 heichips25_sap3/net239 heichips25_sap3/net238 VPWR VGND
+ sg13g2_buf_1
XFILLER_19_880 VPWR VGND sg13g2_decap_4
Xheichips25_sap3_fanout216 heichips25_sap3/net218 heichips25_sap3/net216 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout249 heichips25_sap3/_1451_ heichips25_sap3/net249 VPWR VGND
+ sg13g2_buf_1
Xheichips25_can_lehmann_fsm__1794_ heichips25_can_lehmann_fsm/_1109_ VPWR heichips25_can_lehmann_fsm/_1110_
+ VGND heichips25_can_lehmann_fsm/_0885_ heichips25_can_lehmann_fsm/_0991_ sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2415_ VGND VPWR heichips25_can_lehmann_fsm/_0946_ heichips25_can_lehmann_fsm/net424
+ heichips25_can_lehmann_fsm/_0107_ heichips25_can_lehmann_fsm/_0673_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2346_ heichips25_can_lehmann_fsm/net494 VPWR heichips25_can_lehmann_fsm/_0639_
+ VGND heichips25_can_lehmann_fsm/net1115 heichips25_can_lehmann_fsm/net406 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2277_ heichips25_can_lehmann_fsm/net172 heichips25_can_lehmann_fsm/_0591_
+ heichips25_can_lehmann_fsm/_0592_ VPWR VGND sg13g2_nor2_1
Xheichips25_can_lehmann_fsm_fanout164 heichips25_can_lehmann_fsm/net165 heichips25_can_lehmann_fsm/net164
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout175 heichips25_can_lehmann_fsm/_0495_ heichips25_can_lehmann_fsm/net175
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout186 heichips25_can_lehmann_fsm/net187 heichips25_can_lehmann_fsm/net186
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout197 heichips25_can_lehmann_fsm/net200 heichips25_can_lehmann_fsm/net197
+ VPWR VGND sg13g2_buf_1
XFILLER_0_459 VPWR VGND sg13g2_decap_4
XFILLER_28_110 VPWR VGND sg13g2_fill_1
XFILLER_28_132 VPWR VGND sg13g2_decap_8
XFILLER_17_828 VPWR VGND sg13g2_decap_8
XFILLER_45_55 VPWR VGND sg13g2_fill_2
XFILLER_45_44 VPWR VGND sg13g2_fill_1
XFILLER_43_124 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2160_ heichips25_sap3/_1560_ VPWR heichips25_sap3/_1581_ VGND heichips25_sap3/_1552_
+ heichips25_sap3/_1567_ sg13g2_o21ai_1
XFILLER_45_88 VPWR VGND sg13g2_fill_2
XFILLER_45_66 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2091_ heichips25_sap3/net257 heichips25_sap3/_1438_ heichips25_sap3/net255
+ heichips25_sap3/_1512_ VGND VPWR heichips25_sap3/_1511_ sg13g2_nor4_2
Xheichips25_can_lehmann_fsm__2998__610 VPWR VGND net609 sg13g2_tiehi
XFILLER_12_566 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2993_ heichips25_sap3/_0055_ heichips25_sap3/_0621_ heichips25_sap3/_0622_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__1944_ VPWR heichips25_sap3/_1370_ heichips25_sap3__3998_/Q VGND
+ sg13g2_inv_1
XFILLER_3_231 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3614_ heichips25_sap3/_0876_ heichips25_sap3/_1056_ heichips25_sap3/net140
+ heichips25_sap3/_1179_ VPWR VGND sg13g2_nand3_1
XFILLER_0_971 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3545_ heichips25_sap3/_1134_ heichips25_sap3/_1088_ heichips25_sap3/net144
+ VPWR VGND sg13g2_nand2b_1
XFILLER_47_430 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3476_ VGND VPWR heichips25_sap3/_1411_ heichips25_sap3/net57 heichips25_sap3/_0085_
+ heichips25_sap3/_1075_ sg13g2_a21oi_1
Xheichips25_sap3__2427_ VGND VPWR heichips25_sap3/_1839_ heichips25_sap3/_1843_ heichips25_sap3/_1844_
+ heichips25_sap3/net66 sg13g2_a21oi_1
XFILLER_19_187 VPWR VGND sg13g2_fill_2
XFILLER_34_124 VPWR VGND sg13g2_decap_4
XFILLER_35_658 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2358_ heichips25_sap3/net223 heichips25_sap3/_1777_ heichips25_sap3/_1778_
+ heichips25_sap3/_1779_ VPWR VGND sg13g2_nor3_1
XFILLER_34_157 VPWR VGND sg13g2_decap_4
XFILLER_37_1011 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2289_ heichips25_sap3/_1710_ heichips25_sap3/_1453_ heichips25_sap3/_1709_
+ VPWR VGND sg13g2_nand2_1
XFILLER_34_168 VPWR VGND sg13g2_fill_2
XFILLER_15_382 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__4028_ heichips25_sap3/net458 VGND VPWR heichips25_sap3/net833 heichips25_sap3__4074_/A
+ clknet_leaf_1_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2200_ heichips25_can_lehmann_fsm/_0531_ heichips25_can_lehmann_fsm/net1218
+ heichips25_can_lehmann_fsm/_1101_ VPWR VGND sg13g2_xnor2_1
Xheichips25_can_lehmann_fsm__2131_ heichips25_can_lehmann_fsm/_0470_ heichips25_can_lehmann_fsm/net332
+ heichips25_can_lehmann_fsm__3054_/Q heichips25_can_lehmann_fsm/net319 heichips25_can_lehmann_fsm__3006_/Q
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2062_ heichips25_can_lehmann_fsm/net322 VPWR heichips25_can_lehmann_fsm/_0410_
+ VGND heichips25_can_lehmann_fsm/net179 heichips25_can_lehmann_fsm/_0409_ sg13g2_o21ai_1
XFILLER_38_430 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2964_ net768 VGND VPWR heichips25_can_lehmann_fsm/_0189_
+ heichips25_can_lehmann_fsm__2964_/Q clknet_leaf_18_clk sg13g2_dfrbpq_1
XFILLER_26_603 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1915_ heichips25_can_lehmann_fsm/_1228_ heichips25_can_lehmann_fsm/net333
+ heichips25_can_lehmann_fsm__3051_/Q heichips25_can_lehmann_fsm/net308 heichips25_can_lehmann_fsm__2955_/Q
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2895_ net705 VGND VPWR heichips25_can_lehmann_fsm/net866
+ heichips25_can_lehmann_fsm__2895_/Q clknet_leaf_19_clk sg13g2_dfrbpq_1
X_18__520 VPWR VGND net519 sg13g2_tielo
XFILLER_26_647 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__1846_ heichips25_can_lehmann_fsm/_1152_ heichips25_can_lehmann_fsm/_1142_
+ heichips25_can_lehmann_fsm/_1160_ heichips25_can_lehmann_fsm/_1162_ VPWR VGND sg13g2_a21o_1
Xheichips25_can_lehmann_fsm_hold1114 heichips25_can_lehmann_fsm__2840_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1113 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__1777_ heichips25_can_lehmann_fsm/_1093_ heichips25_can_lehmann_fsm/net305
+ heichips25_can_lehmann_fsm__2941_/Q heichips25_can_lehmann_fsm/net314 heichips25_can_lehmann_fsm__2917_/Q
+ VPWR VGND sg13g2_a22oi_1
XFILLER_15_47 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm_hold1103 heichips25_can_lehmann_fsm__2906_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1102 sg13g2_dlygate4sd3_1
XFILLER_40_127 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm_hold1136 heichips25_can_lehmann_fsm__2916_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1135 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1147 heichips25_can_lehmann_fsm__3021_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1146 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1169 heichips25_can_lehmann_fsm__2833_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1168 sg13g2_dlygate4sd3_1
Xclkbuf_5_5__f_heichips25_sap3\_sap_3_inst.alu_inst.clk heichips25_sap3__3988_/CLK
+ clknet_4_2_0_heichips25_sap3\/sap_3_inst.alu_inst.clk VPWR VGND sg13g2_buf_16
Xheichips25_sap3_hold834 heichips25_sap3/_0169_ VPWR VGND heichips25_sap3/net833 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1158 heichips25_can_lehmann_fsm__3050_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1157 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__2329_ VGND VPWR heichips25_can_lehmann_fsm/_0969_ heichips25_can_lehmann_fsm/net363
+ heichips25_can_lehmann_fsm/_0064_ heichips25_can_lehmann_fsm/_0630_ sg13g2_a21oi_1
Xheichips25_sap3_fanout55 heichips25_sap3/_0748_ heichips25_sap3/net55 VPWR VGND sg13g2_buf_1
Xoutput24 net24 uio_oe[5] VPWR VGND sg13g2_buf_1
Xheichips25_sap3_fanout66 heichips25_sap3/net67 heichips25_sap3/net66 VPWR VGND sg13g2_buf_1
Xheichips25_sap3_fanout77 heichips25_sap3/net78 heichips25_sap3/net77 VPWR VGND sg13g2_buf_1
Xoutput35 net35 uo_out[0] VPWR VGND sg13g2_buf_1
Xheichips25_sap3_fanout88 heichips25_sap3/_1735_ heichips25_sap3/net88 VPWR VGND sg13g2_buf_1
Xheichips25_sap3_fanout99 heichips25_sap3/_0862_ heichips25_sap3/net99 VPWR VGND sg13g2_buf_1
XFILLER_0_267 VPWR VGND sg13g2_fill_1
XFILLER_48_227 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3330_ heichips25_sap3/_0940_ heichips25_sap3/net138 heichips25_sap3__3974_/Q
+ heichips25_sap3/net140 heichips25_sap3__3982_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3261_ VGND VPWR heichips25_sap3/net59 heichips25_sap3/_0870_ heichips25_sap3/_0874_
+ heichips25_sap3/_0777_ sg13g2_a21oi_1
Xheichips25_sap3__2212_ heichips25_sap3/_1578_ heichips25_sap3/_1617_ heichips25_sap3/_1628_
+ heichips25_sap3/_1632_ heichips25_sap3/_1633_ VPWR VGND sg13g2_nor4_1
XFILLER_16_102 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3192_ heichips25_sap3/_0805_ heichips25_sap3__4007_/Q heichips25_sap3/net148
+ VPWR VGND sg13g2_nand2_1
XFILLER_32_606 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2143_ VPWR VGND heichips25_sap3/_1522_ heichips25_sap3/_1562_ heichips25_sap3/_1563_
+ heichips25_sap3/_1524_ heichips25_sap3/_1564_ heichips25_sap3/_1534_ sg13g2_a221oi_1
XFILLER_16_168 VPWR VGND sg13g2_fill_2
XFILLER_32_628 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2074_ heichips25_sap3/_1487_ heichips25_sap3/_1489_ heichips25_sap3/_1436_
+ heichips25_sap3/_1495_ VPWR VGND sg13g2_nand3_1
Xheichips25_sap3_hold1180 heichips25_sap3/_0182_ VPWR VGND heichips25_sap3/net1179
+ sg13g2_dlygate4sd3_1
XFILLER_8_334 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2902__692 VPWR VGND net691 sg13g2_tiehi
XFILLER_4_551 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2976_ heichips25_sap3/_0049_ heichips25_sap3/_0610_ heichips25_sap3/_0611_
+ VPWR VGND sg13g2_nand2_1
XFILLER_39_205 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3528_ heichips25_sap3/_1116_ heichips25_sap3/_1119_ heichips25_sap3/_1120_
+ VPWR VGND sg13g2_nor2_1
XFILLER_11_4 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1700_ heichips25_can_lehmann_fsm/_1024_ heichips25_can_lehmann_fsm/net296
+ heichips25_can_lehmann_fsm__2895_/Q heichips25_can_lehmann_fsm/net313 heichips25_can_lehmann_fsm__2919_/Q
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3459_ heichips25_sap3/_1061_ heichips25_sap3/_1062_ heichips25_sap3/_1063_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_can_lehmann_fsm__2680_ heichips25_can_lehmann_fsm/net464 VPWR heichips25_can_lehmann_fsm/_0806_
+ VGND heichips25_can_lehmann_fsm/net924 heichips25_can_lehmann_fsm/net357 sg13g2_o21ai_1
XFILLER_35_488 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1631_ VPWR heichips25_can_lehmann_fsm/_0955_ heichips25_can_lehmann_fsm/net922
+ VGND sg13g2_inv_1
XFILLER_22_138 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__1562_ VPWR heichips25_can_lehmann_fsm/_0886_ heichips25_can_lehmann_fsm/net1090
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__2114_ VGND VPWR heichips25_can_lehmann_fsm/_0943_ heichips25_can_lehmann_fsm/net303
+ heichips25_can_lehmann_fsm/_0453_ heichips25_can_lehmann_fsm/_0452_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2834__539 VPWR VGND net538 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2045_ VPWR VGND heichips25_can_lehmann_fsm/_0392_ heichips25_can_lehmann_fsm/net193
+ heichips25_can_lehmann_fsm/net189 heichips25_can_lehmann_fsm__2791_/Q heichips25_can_lehmann_fsm/_0394_
+ heichips25_can_lehmann_fsm/net198 sg13g2_a221oi_1
Xheichips25_can_lehmann_fsm__2947_ net547 VGND VPWR heichips25_can_lehmann_fsm/net935
+ heichips25_can_lehmann_fsm__2947_/Q clknet_leaf_21_clk sg13g2_dfrbpq_1
XFILLER_38_293 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2878_ net739 VGND VPWR heichips25_can_lehmann_fsm/_0103_
+ heichips25_can_lehmann_fsm__2878_/Q clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_13_105 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1829_ heichips25_can_lehmann_fsm/_1145_ heichips25_can_lehmann_fsm/net343
+ net6 VPWR VGND sg13g2_nand2_1
XFILLER_26_499 VPWR VGND sg13g2_decap_4
XFILLER_42_959 VPWR VGND sg13g2_fill_1
XFILLER_13_138 VPWR VGND sg13g2_decap_4
XFILLER_10_801 VPWR VGND sg13g2_fill_2
XFILLER_22_650 VPWR VGND sg13g2_decap_4
XFILLER_42_78 VPWR VGND sg13g2_decap_4
XFILLER_6_838 VPWR VGND sg13g2_fill_2
XFILLER_5_315 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2830_ VGND VPWR heichips25_sap3__3908_/Q heichips25_sap3/net204
+ heichips25_sap3/_0474_ heichips25_sap3/net158 sg13g2_a21oi_1
Xheichips25_sap3__2761_ heichips25_sap3/_0406_ heichips25_sap3/_0405_ heichips25_sap3/_0407_
+ VPWR VGND sg13g2_nor2b_1
Xheichips25_sap3__2692_ heichips25_sap3/_1887_ heichips25_sap3/_0337_ heichips25_sap3/_0338_
+ VPWR VGND sg13g2_nor2_1
XFILLER_3_28 VPWR VGND sg13g2_decap_8
XFILLER_49_525 VPWR VGND sg13g2_decap_8
XFILLER_49_569 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3313_ heichips25_sap3/net119 heichips25_sap3/_0923_ heichips25_sap3/_0924_
+ VPWR VGND sg13g2_nor2_1
XFILLER_17_422 VPWR VGND sg13g2_decap_8
XFILLER_29_260 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3244_ heichips25_sap3/_0795_ heichips25_sap3/_0802_ heichips25_sap3/net63
+ heichips25_sap3/_0855_ heichips25_sap3/_0857_ VPWR VGND sg13g2_nor4_1
XFILLER_33_904 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3175_ heichips25_sap3/_0788_ heichips25_sap3/net135 heichips25_sap3__3977_/Q
+ heichips25_sap3/net142 heichips25_sap3__3993_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2126_ heichips25_sap3/_1547_ heichips25_sap3/net250 heichips25_sap3/net251
+ VPWR VGND sg13g2_nand2b_1
XFILLER_9_621 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2057_ heichips25_sap3/_1478_ heichips25_sap3/net251 heichips25_sap3/net250
+ VPWR VGND sg13g2_nand2b_1
XFILLER_9_676 VPWR VGND sg13g2_fill_1
XFILLER_8_175 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2959_ heichips25_sap3/_0592_ heichips25_sap3/_0595_ heichips25_sap3/_0591_
+ heichips25_sap3/_0597_ VPWR VGND heichips25_sap3/_0596_ sg13g2_nand4_1
Xheichips25_can_lehmann_fsm__2801_ net604 VGND VPWR heichips25_can_lehmann_fsm/_0026_
+ heichips25_can_lehmann_fsm__2801_/Q clknet_leaf_4_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2732_ heichips25_can_lehmann_fsm/net466 VPWR heichips25_can_lehmann_fsm/_0832_
+ VGND heichips25_can_lehmann_fsm/net908 heichips25_can_lehmann_fsm/net393 sg13g2_o21ai_1
XFILLER_24_904 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2663_ VGND VPWR heichips25_can_lehmann_fsm/_0880_ heichips25_can_lehmann_fsm/net418
+ heichips25_can_lehmann_fsm/_0231_ heichips25_can_lehmann_fsm/_0797_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__1614_ VPWR heichips25_can_lehmann_fsm/_0938_ heichips25_can_lehmann_fsm/net1100
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__2594_ heichips25_can_lehmann_fsm/net480 VPWR heichips25_can_lehmann_fsm/_0763_
+ VGND heichips25_can_lehmann_fsm/net972 heichips25_can_lehmann_fsm/net399 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__1545_ VPWR heichips25_can_lehmann_fsm/_0869_ heichips25_can_lehmann_fsm/net960
+ VGND sg13g2_inv_1
XFILLER_31_480 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2028_ VGND VPWR heichips25_can_lehmann_fsm/net1238 heichips25_can_lehmann_fsm/net189
+ heichips25_can_lehmann_fsm/_0379_ heichips25_can_lehmann_fsm/net193 sg13g2_a21oi_1
XFILLER_46_517 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2886__724 VPWR VGND net723 sg13g2_tiehi
XFILLER_37_78 VPWR VGND sg13g2_fill_1
XFILLER_42_723 VPWR VGND sg13g2_fill_2
XFILLER_14_403 VPWR VGND sg13g2_decap_8
XFILLER_15_926 VPWR VGND sg13g2_fill_1
XFILLER_41_266 VPWR VGND sg13g2_fill_2
XFILLER_23_992 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3931_ heichips25_sap3/net438 VGND VPWR heichips25_sap3/_0072_ heichips25_sap3__3931_/Q
+ clkload18/A sg13g2_dfrbpq_1
XFILLER_5_145 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3862_ heichips25_sap3/_1357_ VPWR heichips25_sap3/_0189_ VGND heichips25_sap3/_1359_
+ heichips25_sap3/_1433_ sg13g2_o21ai_1
XFILLER_5_189 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2813_ heichips25_sap3/net70 heichips25_sap3/net289 heichips25_sap3/_0457_
+ heichips25_sap3/_0040_ VPWR VGND sg13g2_a21o_1
Xheichips25_sap3__3793_ heichips25_sap3/net339 heichips25_sap3/net1120 heichips25_sap3/_1302_
+ heichips25_sap3/_0175_ VPWR VGND sg13g2_a21o_1
Xheichips25_sap3__2744_ heichips25_sap3/_0363_ heichips25_sap3/_0389_ heichips25_sap3/_0390_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__2675_ heichips25_sap3/net288 heichips25_sap3__3882_/Q heichips25_sap3/_0297_
+ heichips25_sap3/_0023_ VPWR VGND sg13g2_mux2_1
Xclkbuf_5_23__f_heichips25_sap3\_sap_3_inst.alu_inst.clk clkload26/A clknet_4_11_0_heichips25_sap3\/sap_3_inst.alu_inst.clk
+ VPWR VGND sg13g2_buf_16
XFILLER_37_517 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2787__633 VPWR VGND net632 sg13g2_tiehi
XFILLER_17_263 VPWR VGND sg13g2_decap_8
XFILLER_45_594 VPWR VGND sg13g2_fill_1
XFILLER_45_583 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3227_ heichips25_sap3/_0836_ heichips25_sap3/_0837_ heichips25_sap3/_0838_
+ heichips25_sap3/_0839_ heichips25_sap3/_0840_ VPWR VGND sg13g2_and4_1
XFILLER_32_211 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3158_ heichips25_sap3/_0771_ heichips25_sap3/_0680_ heichips25_sap3/_0696_
+ VPWR VGND sg13g2_nand2_1
XFILLER_32_233 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2109_ heichips25_sap3/net267 heichips25_sap3/_1529_ heichips25_sap3/_1530_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__3089_ heichips25_sap3/_0702_ heichips25_sap3/_1560_ heichips25_sap3/net222
+ VPWR VGND sg13g2_nand2_1
XFILLER_14_992 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__3000_ net593 VGND VPWR heichips25_can_lehmann_fsm/net845
+ heichips25_can_lehmann_fsm__3000_/Q clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_4_60 VPWR VGND sg13g2_decap_8
XFILLER_43_509 VPWR VGND sg13g2_decap_8
XFILLER_36_550 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2715_ VGND VPWR heichips25_can_lehmann_fsm/_0866_ heichips25_can_lehmann_fsm/net378
+ heichips25_can_lehmann_fsm/_0257_ heichips25_can_lehmann_fsm/_0823_ sg13g2_a21oi_1
XFILLER_23_233 VPWR VGND sg13g2_fill_2
XFILLER_23_244 VPWR VGND sg13g2_decap_8
XFILLER_24_789 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2646_ heichips25_can_lehmann_fsm/net472 VPWR heichips25_can_lehmann_fsm/_0789_
+ VGND heichips25_can_lehmann_fsm__2998_/Q heichips25_can_lehmann_fsm/net404 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2577_ VGND VPWR heichips25_can_lehmann_fsm/_0903_ heichips25_can_lehmann_fsm/net370
+ heichips25_can_lehmann_fsm/_0188_ heichips25_can_lehmann_fsm/_0754_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__1528_ VPWR heichips25_can_lehmann_fsm/_0852_ heichips25_can_lehmann_fsm/net1132
+ VGND sg13g2_inv_1
Xheichips25_sap3__2460_ VGND VPWR heichips25_sap3/_1479_ heichips25_sap3/_1623_ heichips25_sap3/_1873_
+ heichips25_sap3/_1872_ sg13g2_a21oi_1
Xheichips25_sap3__2391_ heichips25_sap3/_1804_ heichips25_sap3/_1805_ heichips25_sap3/_1734_
+ heichips25_sap3/_1810_ VPWR VGND heichips25_sap3/_1809_ sg13g2_nand4_1
XFILLER_46_358 VPWR VGND sg13g2_fill_1
XFILLER_0_29 VPWR VGND sg13g2_decap_8
XFILLER_27_550 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__4061_ heichips25_sap3/net459 VGND VPWR heichips25_sap3/_0000_ heichips25_sap3__4061_/Q
+ clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_14_211 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3012_ heichips25_sap3/_0632_ heichips25_sap3/net270 heichips25_sap3/net231
+ VPWR VGND sg13g2_nand2_1
XFILLER_9_38 VPWR VGND sg13g2_decap_8
XFILLER_6_443 VPWR VGND sg13g2_fill_2
XFILLER_10_494 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3914_ heichips25_sap3/net455 VGND VPWR heichips25_sap3/_0055_ heichips25_sap3__3914_/Q
+ clkload26/A sg13g2_dfrbpq_1
Xheichips25_sap3__3845_ heichips25_sap3/_1345_ VPWR heichips25_sap3/_0184_ VGND heichips25_sap3/_0018_
+ heichips25_sap3/_1262_ sg13g2_o21ai_1
Xheichips25_sap3__3776_ heichips25_sap3/_1287_ heichips25_sap3/_1278_ heichips25_sap3__4004_/Q
+ heichips25_sap3/_1259_ heichips25_sap3__3980_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_36_6 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2727_ heichips25_sap3/_0373_ heichips25_sap3/net254 heichips25_sap3/_0372_
+ VPWR VGND sg13g2_nand2_1
XFILLER_49_130 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2658_ VGND VPWR heichips25_sap3/_1679_ heichips25_sap3/_0323_ heichips25_sap3/_0003_
+ heichips25_sap3__4063_/Q sg13g2_a21oi_1
XFILLER_37_314 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2589_ heichips25_sap3/_0262_ heichips25_sap3/net76 heichips25_sap3__3989_/Q
+ heichips25_sap3/net82 heichips25_sap3__3973_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2500_ heichips25_can_lehmann_fsm/net469 VPWR heichips25_can_lehmann_fsm/_0716_
+ VGND heichips25_can_lehmann_fsm/net1054 heichips25_can_lehmann_fsm/net359 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2431_ VGND VPWR heichips25_can_lehmann_fsm/_0940_ heichips25_can_lehmann_fsm/net412
+ heichips25_can_lehmann_fsm/_0115_ heichips25_can_lehmann_fsm/_0681_ sg13g2_a21oi_1
XFILLER_33_575 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2362_ heichips25_can_lehmann_fsm/net500 VPWR heichips25_can_lehmann_fsm/_0647_
+ VGND heichips25_can_lehmann_fsm/net941 heichips25_can_lehmann_fsm/net430 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2293_ VGND VPWR heichips25_can_lehmann_fsm/net948 heichips25_can_lehmann_fsm/net171
+ heichips25_can_lehmann_fsm/_0605_ heichips25_can_lehmann_fsm/_0604_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm_fanout302 heichips25_can_lehmann_fsm/net304 heichips25_can_lehmann_fsm/net302
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout313 heichips25_can_lehmann_fsm/net316 heichips25_can_lehmann_fsm/net313
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout346 heichips25_can_lehmann_fsm/net1219 heichips25_can_lehmann_fsm/net346
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout324 heichips25_can_lehmann_fsm/net330 heichips25_can_lehmann_fsm/net324
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout357 heichips25_can_lehmann_fsm/net358 heichips25_can_lehmann_fsm/net357
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout335 heichips25_can_lehmann_fsm/net336 heichips25_can_lehmann_fsm/net335
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout368 heichips25_can_lehmann_fsm/net369 heichips25_can_lehmann_fsm/net368
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout379 heichips25_can_lehmann_fsm/net389 heichips25_can_lehmann_fsm/net379
+ VPWR VGND sg13g2_buf_1
XFILLER_29_848 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2963__773 VPWR VGND net772 sg13g2_tiehi
XFILLER_24_531 VPWR VGND sg13g2_decap_8
XFILLER_24_553 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2629_ VGND VPWR heichips25_can_lehmann_fsm/_0890_ heichips25_can_lehmann_fsm/net368
+ heichips25_can_lehmann_fsm/_0214_ heichips25_can_lehmann_fsm/_0780_ sg13g2_a21oi_1
XFILLER_12_715 VPWR VGND sg13g2_fill_1
XFILLER_11_247 VPWR VGND sg13g2_fill_2
XFILLER_12_748 VPWR VGND sg13g2_fill_2
XFILLER_7_207 VPWR VGND sg13g2_decap_8
Xclkload1 clkload1/Y clknet_leaf_1_clk VPWR VGND sg13g2_inv_2
Xheichips25_sap3__1960_ VPWR heichips25_sap3/_1386_ heichips25_sap3__4012_/Q VGND
+ sg13g2_inv_1
Xheichips25_sap3__3630_ VGND VPWR heichips25_sap3/net142 heichips25_sap3/_0881_ heichips25_sap3/_1187_
+ heichips25_sap3/net132 sg13g2_a21oi_1
Xheichips25_sap3__3561_ heichips25_sap3/_1142_ heichips25_sap3__3963_/Q heichips25_sap3/net100
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__2512_ heichips25_sap3/_1899_ VPWR heichips25_sap3/_1924_ VGND heichips25_sap3/_1802_
+ uio_out_sap3\[1\] sg13g2_o21ai_1
Xheichips25_sap3__3492_ uio_oe_sap3\[0\] heichips25_sap3/_1088_ heichips25_sap3/_1089_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__2443_ heichips25_sap3/_1858_ heichips25_sap3/net73 heichips25_sap3__4007_/Q
+ heichips25_sap3/net81 heichips25_sap3__3975_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2374_ heichips25_sap3/_1793_ heichips25_sap3/_1794_ heichips25_sap3/_1795_
+ VPWR VGND sg13g2_and2_1
XFILLER_15_520 VPWR VGND sg13g2_decap_8
XFILLER_28_881 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__4044_ heichips25_sap3/net452 VGND VPWR heichips25_sap3/net839 heichips25_sap3__4071_/A
+ clknet_leaf_22_clk sg13g2_dfrbpq_1
XFILLER_42_350 VPWR VGND sg13g2_decap_4
XFILLER_30_512 VPWR VGND sg13g2_decap_8
XFILLER_30_523 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_hold980 heichips25_can_lehmann_fsm/_0211_ VPWR VGND heichips25_can_lehmann_fsm/net979
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold991 heichips25_can_lehmann_fsm__3019_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net990 sg13g2_dlygate4sd3_1
Xheichips25_sap3__3828_ VPWR VGND heichips25_sap3/_1333_ heichips25_sap3/net340 heichips25_sap3/_1328_
+ heichips25_sap3/_1412_ heichips25_sap3/_1334_ heichips25_sap3/net291 sg13g2_a221oi_1
Xheichips25_sap3__3759_ heichips25_sap3/_1271_ heichips25_sap3__4040_/Q heichips25_sap3__4041_/Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_3_991 VPWR VGND sg13g2_decap_8
XFILLER_2_490 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2980_ net704 VGND VPWR heichips25_can_lehmann_fsm/net873
+ heichips25_can_lehmann_fsm__2980_/Q clknet_leaf_14_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1931_ VGND VPWR heichips25_can_lehmann_fsm__3050_/Q heichips25_can_lehmann_fsm/_1161_
+ heichips25_can_lehmann_fsm/_0294_ heichips25_can_lehmann_fsm/_1139_ sg13g2_a21oi_1
XFILLER_37_133 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2912__672 VPWR VGND net671 sg13g2_tiehi
X_27_ net512 net829 net506 net24 VPWR VGND sg13g2_mux2_1
Xheichips25_can_lehmann_fsm__1862_ heichips25_can_lehmann_fsm/_1176_ heichips25_can_lehmann_fsm/_1177_
+ heichips25_can_lehmann_fsm/_0000_ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3_fanout217 heichips25_sap3/net218 heichips25_sap3/net217 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout228 heichips25_sap3/_1597_ heichips25_sap3/net228 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout239 heichips25_sap3/net240 heichips25_sap3/net239 VPWR VGND
+ sg13g2_buf_1
Xheichips25_can_lehmann_fsm__1793_ heichips25_can_lehmann_fsm/net350 heichips25_can_lehmann_fsm/net351
+ heichips25_can_lehmann_fsm__3045_/Q heichips25_can_lehmann_fsm/_1109_ VPWR VGND
+ heichips25_can_lehmann_fsm/net354 sg13g2_nand4_1
XFILLER_40_309 VPWR VGND sg13g2_fill_1
XFILLER_33_361 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2414_ heichips25_can_lehmann_fsm/net500 VPWR heichips25_can_lehmann_fsm/_0673_
+ VGND heichips25_can_lehmann_fsm/net879 heichips25_can_lehmann_fsm/net430 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2345_ VGND VPWR heichips25_can_lehmann_fsm/_0965_ heichips25_can_lehmann_fsm/net367
+ heichips25_can_lehmann_fsm/_0072_ heichips25_can_lehmann_fsm/_0638_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2276_ heichips25_can_lehmann_fsm/_1047_ heichips25_can_lehmann_fsm/net1191
+ heichips25_can_lehmann_fsm/_0591_ VPWR VGND sg13g2_xor2_1
Xheichips25_can_lehmann_fsm_fanout165 heichips25_can_lehmann_fsm/_0496_ heichips25_can_lehmann_fsm/net165
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout176 heichips25_can_lehmann_fsm/_0495_ heichips25_can_lehmann_fsm/net176
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout187 heichips25_can_lehmann_fsm/_0309_ heichips25_can_lehmann_fsm/net187
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout198 heichips25_can_lehmann_fsm/net200 heichips25_can_lehmann_fsm/net198
+ VPWR VGND sg13g2_buf_1
XFILLER_29_79 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2813__581 VPWR VGND net580 sg13g2_tiehi
XFILLER_28_177 VPWR VGND sg13g2_decap_8
XFILLER_28_188 VPWR VGND sg13g2_fill_2
XFILLER_28_199 VPWR VGND sg13g2_decap_8
XFILLER_43_169 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2090_ heichips25_sap3/net266 heichips25_sap3/net272 heichips25_sap3/_1511_
+ VPWR VGND heichips25_sap3/net269 sg13g2_nand3b_1
XFILLER_24_372 VPWR VGND sg13g2_fill_1
XFILLER_31_309 VPWR VGND sg13g2_decap_4
XFILLER_12_534 VPWR VGND sg13g2_decap_8
XFILLER_8_538 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2992_ heichips25_sap3/_0622_ heichips25_sap3/_0606_ heichips25_sap3/_0412_
+ heichips25_sap3/_0605_ heichips25_sap3/net275 VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__1943_ VPWR heichips25_sap3/_1369_ heichips25_sap3__4014_/Q VGND
+ sg13g2_inv_1
XFILLER_3_254 VPWR VGND sg13g2_fill_2
XFILLER_3_243 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3613_ heichips25_sap3/_1178_ VPWR heichips25_sap3/_0119_ VGND heichips25_sap3/_1171_
+ heichips25_sap3/_1177_ sg13g2_o21ai_1
XFILLER_3_287 VPWR VGND sg13g2_decap_8
XFILLER_10_81 VPWR VGND sg13g2_decap_8
XFILLER_0_950 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3544_ heichips25_sap3/_0095_ heichips25_sap3/_1130_ heichips25_sap3/_1133_
+ heichips25_sap3/net107 heichips25_sap3/_1425_ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3475_ heichips25_sap3/net57 heichips25_sap3/_1073_ heichips25_sap3/_1074_
+ heichips25_sap3/_1075_ VPWR VGND sg13g2_nor3_1
Xheichips25_sap3__2426_ heichips25_sap3/_1843_ heichips25_sap3/_1840_ heichips25_sap3/_1841_
+ heichips25_sap3/_1842_ VPWR VGND sg13g2_and3_1
XFILLER_37_1001 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2357_ VGND VPWR heichips25_sap3/net229 heichips25_sap3/_1550_ heichips25_sap3/_1778_
+ heichips25_sap3/_1518_ sg13g2_a21oi_1
XFILLER_16_851 VPWR VGND sg13g2_fill_1
XFILLER_34_147 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2288_ heichips25_sap3/_1709_ heichips25_sap3/net270 heichips25_sap3/_1651_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__4027_ heichips25_sap3/net461 VGND VPWR heichips25_sap3/net1059 heichips25_sap3__4073_/A
+ clknet_leaf_2_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2977__717 VPWR VGND net716 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2130_ heichips25_can_lehmann_fsm/net337 VPWR heichips25_can_lehmann_fsm/_0469_
+ VGND heichips25_can_lehmann_fsm__2982_/Q heichips25_can_lehmann_fsm/_0983_ sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2061_ heichips25_can_lehmann_fsm/_0409_ heichips25_can_lehmann_fsm/_0304_
+ heichips25_can_lehmann_fsm__2793_/Q VPWR VGND sg13g2_nand2b_1
Xheichips25_can_lehmann_fsm__2963_ net772 VGND VPWR heichips25_can_lehmann_fsm/_0188_
+ heichips25_can_lehmann_fsm__2963_/Q clknet_leaf_18_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2894_ net707 VGND VPWR heichips25_can_lehmann_fsm/net1101
+ heichips25_can_lehmann_fsm__2894_/Q clknet_leaf_19_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1914_ heichips25_can_lehmann_fsm/_1227_ heichips25_can_lehmann_fsm/_1226_
+ heichips25_can_lehmann_fsm/net337 heichips25_can_lehmann_fsm/net297 heichips25_can_lehmann_fsm__2907_/Q
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__1845_ VPWR VGND heichips25_can_lehmann_fsm__3060_/Q heichips25_can_lehmann_fsm/_1159_
+ heichips25_can_lehmann_fsm/_1153_ heichips25_can_lehmann_fsm/_1142_ heichips25_can_lehmann_fsm/_1161_
+ heichips25_can_lehmann_fsm/_1152_ sg13g2_a221oi_1
Xheichips25_can_lehmann_fsm__2845__806 VPWR VGND net805 sg13g2_tiehi
XFILLER_25_125 VPWR VGND sg13g2_fill_1
XFILLER_26_659 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_hold1115 heichips25_can_lehmann_fsm__3023_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1114 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1104 heichips25_can_lehmann_fsm__2953_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1103 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__1776_ heichips25_can_lehmann_fsm/_1092_ heichips25_can_lehmann_fsm/net295
+ heichips25_can_lehmann_fsm__2965_/Q heichips25_can_lehmann_fsm/net296 heichips25_can_lehmann_fsm__2893_/Q
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm_hold1137 heichips25_can_lehmann_fsm__2836_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1136 sg13g2_dlygate4sd3_1
XFILLER_21_320 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_hold1148 heichips25_can_lehmann_fsm__3047_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1147 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1159 heichips25_can_lehmann_fsm__2831_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1158 sg13g2_dlygate4sd3_1
XFILLER_22_876 VPWR VGND sg13g2_fill_2
XFILLER_21_375 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2328_ heichips25_can_lehmann_fsm/net471 VPWR heichips25_can_lehmann_fsm/_0630_
+ VGND heichips25_can_lehmann_fsm/net933 heichips25_can_lehmann_fsm/net363 sg13g2_o21ai_1
Xheichips25_sap3_fanout45 heichips25_sap3/_0242_ heichips25_sap3/net45 VPWR VGND sg13g2_buf_2
Xheichips25_can_lehmann_fsm__2259_ VGND VPWR heichips25_can_lehmann_fsm/net206 heichips25_can_lehmann_fsm/net1184
+ heichips25_can_lehmann_fsm/_0047_ heichips25_can_lehmann_fsm/_0577_ sg13g2_a21oi_1
Xheichips25_sap3_fanout67 heichips25_sap3/_1593_ heichips25_sap3/net67 VPWR VGND sg13g2_buf_1
Xheichips25_sap3_fanout78 heichips25_sap3/_1743_ heichips25_sap3/net78 VPWR VGND sg13g2_buf_1
Xheichips25_sap3_fanout56 heichips25_sap3/_1134_ heichips25_sap3/net56 VPWR VGND sg13g2_buf_1
Xoutput25 net25 uio_oe[6] VPWR VGND sg13g2_buf_1
Xoutput36 net36 uo_out[1] VPWR VGND sg13g2_buf_1
Xheichips25_sap3_fanout89 heichips25_sap3/net92 heichips25_sap3/net89 VPWR VGND sg13g2_buf_1
XFILLER_0_246 VPWR VGND sg13g2_decap_8
XFILLER_0_213 VPWR VGND sg13g2_decap_8
XFILLER_5_1010 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3260_ heichips25_sap3/_0794_ heichips25_sap3/net61 heichips25_sap3/_0868_
+ heichips25_sap3/_0873_ VPWR VGND sg13g2_nor3_1
Xheichips25_sap3__2211_ heichips25_sap3/_1448_ heichips25_sap3/net234 heichips25_sap3/_1488_
+ heichips25_sap3/_1632_ VPWR VGND sg13g2_nor3_1
XFILLER_17_615 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3191_ heichips25_sap3/_0804_ heichips25_sap3/net132 heichips25_sap3__3999_/Q
+ heichips25_sap3/net135 heichips25_sap3__3975_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2142_ heichips25_sap3/_1563_ heichips25_sap3/_1498_ heichips25_sap3/_1560_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__2073_ heichips25_sap3/_1437_ heichips25_sap3/net255 heichips25_sap3/_1490_
+ heichips25_sap3/_1494_ VPWR VGND sg13g2_nor3_1
XFILLER_25_692 VPWR VGND sg13g2_fill_1
XFILLER_9_803 VPWR VGND sg13g2_decap_8
XFILLER_12_331 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2896__704 VPWR VGND net703 sg13g2_tiehi
XFILLER_12_375 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2975_ heichips25_sap3/_0611_ heichips25_sap3/net153 heichips25_sap3/_0400_
+ heichips25_sap3/net167 heichips25_sap3/net286 VPWR VGND sg13g2_a22oi_1
XFILLER_39_239 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3527_ heichips25_sap3/net109 VPWR heichips25_sap3/_1119_ VGND heichips25_sap3/_1117_
+ heichips25_sap3/_1118_ sg13g2_o21ai_1
XFILLER_0_791 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3458_ heichips25_sap3/_0863_ heichips25_sap3/_0903_ heichips25_sap3/_1062_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__2409_ heichips25_sap3/_1826_ heichips25_sap3/net75 heichips25_sap3__3984_/Q
+ heichips25_sap3/net81 heichips25_sap3__3968_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3389_ heichips25_sap3/_0996_ VPWR heichips25_sap3/_0997_ VGND heichips25_sap3/net123
+ heichips25_sap3/_0994_ sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__1630_ VPWR heichips25_can_lehmann_fsm/_0954_ heichips25_can_lehmann_fsm/net987
+ VGND sg13g2_inv_1
XFILLER_22_106 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1561_ VPWR heichips25_can_lehmann_fsm/_0885_ heichips25_can_lehmann_fsm/net855
+ VGND sg13g2_inv_1
XFILLER_15_191 VPWR VGND sg13g2_decap_4
XFILLER_30_161 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2797__613 VPWR VGND net612 sg13g2_tiehi
XFILLER_30_183 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2113_ VPWR VGND heichips25_can_lehmann_fsm__3053_/Q heichips25_can_lehmann_fsm/_0451_
+ heichips25_can_lehmann_fsm/net333 heichips25_can_lehmann_fsm__3005_/Q heichips25_can_lehmann_fsm/_0452_
+ heichips25_can_lehmann_fsm/net319 sg13g2_a221oi_1
Xheichips25_can_lehmann_fsm__2044_ heichips25_can_lehmann_fsm/_0982_ heichips25_can_lehmann_fsm/net193
+ heichips25_can_lehmann_fsm/_0393_ VPWR VGND sg13g2_and2_1
Xheichips25_can_lehmann_fsm__2946_ net551 VGND VPWR heichips25_can_lehmann_fsm/net905
+ heichips25_can_lehmann_fsm__2946_/Q clknet_leaf_21_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2877_ net741 VGND VPWR heichips25_can_lehmann_fsm/_0102_
+ heichips25_can_lehmann_fsm__2877_/Q clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_41_415 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1828_ heichips25_can_lehmann_fsm/_1144_ heichips25_can_lehmann_fsm__3044_/Q
+ heichips25_can_lehmann_fsm/_1143_ VPWR VGND sg13g2_nand2_1
Xheichips25_can_lehmann_fsm__1759_ heichips25_can_lehmann_fsm/_1078_ heichips25_can_lehmann_fsm__2790_/Q
+ heichips25_can_lehmann_fsm/_1037_ VPWR VGND sg13g2_nand2_1
XFILLER_42_46 VPWR VGND sg13g2_fill_1
XFILLER_1_511 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2760_ heichips25_sap3/_0406_ heichips25_sap3/_0356_ heichips25_sap3/_0394_
+ VPWR VGND sg13g2_xnor2_1
Xheichips25_sap3__2691_ heichips25_sap3/_0337_ heichips25_sap3/_1884_ heichips25_sap3/net168
+ VPWR VGND sg13g2_nand2_1
XFILLER_49_548 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3312_ heichips25_sap3/net50 heichips25_sap3/_0900_ heichips25_sap3/_0923_
+ VPWR VGND sg13g2_xor2_1
XFILLER_45_743 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3243_ heichips25_sap3/_0802_ heichips25_sap3/net63 heichips25_sap3/_0855_
+ heichips25_sap3/_0856_ VPWR VGND sg13g2_nor3_1
XFILLER_18_968 VPWR VGND sg13g2_fill_1
XFILLER_45_776 VPWR VGND sg13g2_decap_8
XFILLER_44_253 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3174_ heichips25_sap3/_0787_ heichips25_sap3/net132 heichips25_sap3__4001_/Q
+ heichips25_sap3/net139 heichips25_sap3__3985_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_17_478 VPWR VGND sg13g2_decap_8
XFILLER_32_404 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2125_ heichips25_sap3/net251 heichips25_sap3__4066_/Q heichips25_sap3/_1546_
+ VPWR VGND sg13g2_nor2b_1
XFILLER_33_949 VPWR VGND sg13g2_fill_1
XFILLER_41_982 VPWR VGND sg13g2_fill_1
XFILLER_8_121 VPWR VGND sg13g2_fill_1
XFILLER_8_110 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2056_ heichips25_sap3/net250 heichips25_sap3/net251 heichips25_sap3/_1477_
+ VPWR VGND sg13g2_nor2b_1
XFILLER_9_688 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2958_ VGND VPWR heichips25_sap3/_0343_ heichips25_sap3/_0412_ heichips25_sap3/_0596_
+ heichips25_sap3/net65 sg13g2_a21oi_1
XFILLER_5_861 VPWR VGND sg13g2_fill_2
XFILLER_4_393 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2889_ heichips25_sap3/_0530_ heichips25_sap3/net281 heichips25_sap3/net211
+ VPWR VGND sg13g2_xnor2_1
Xheichips25_can_lehmann_fsm__2800_ net606 VGND VPWR heichips25_can_lehmann_fsm/net1271
+ heichips25_can_lehmann_fsm__2800_/Q clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_36_732 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2731_ VGND VPWR heichips25_can_lehmann_fsm/_0862_ heichips25_can_lehmann_fsm/net356
+ heichips25_can_lehmann_fsm/_0265_ heichips25_can_lehmann_fsm/_0831_ sg13g2_a21oi_1
XFILLER_35_242 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2662_ heichips25_can_lehmann_fsm/net488 VPWR heichips25_can_lehmann_fsm/_0797_
+ VGND heichips25_can_lehmann_fsm__3006_/Q heichips25_can_lehmann_fsm/net418 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__1613_ VPWR heichips25_can_lehmann_fsm/_0937_ heichips25_can_lehmann_fsm/net865
+ VGND sg13g2_inv_1
XFILLER_23_448 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2593_ VGND VPWR heichips25_can_lehmann_fsm/_0899_ heichips25_can_lehmann_fsm/net360
+ heichips25_can_lehmann_fsm/_0196_ heichips25_can_lehmann_fsm/_0762_ sg13g2_a21oi_1
XFILLER_23_459 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1544_ VPWR heichips25_can_lehmann_fsm/_0868_ heichips25_can_lehmann_fsm/net1152
+ VGND sg13g2_inv_1
XFILLER_31_470 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2027_ VPWR VGND heichips25_can_lehmann_fsm/net192 heichips25_can_lehmann_fsm/_0378_
+ heichips25_can_lehmann_fsm/_0377_ heichips25_can_lehmann_fsm/_0375_ heichips25_can_lehmann_fsm/_0014_
+ heichips25_can_lehmann_fsm/_0376_ sg13g2_a221oi_1
XFILLER_39_592 VPWR VGND sg13g2_fill_1
XFILLER_26_231 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2929_ net619 VGND VPWR heichips25_can_lehmann_fsm/net859
+ heichips25_can_lehmann_fsm__2929_/Q clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_26_253 VPWR VGND sg13g2_fill_2
Xclkbuf_5_6__f_heichips25_sap3\_sap_3_inst.alu_inst.clk heichips25_sap3__4015_/CLK
+ clknet_4_3_0_heichips25_sap3\/sap_3_inst.alu_inst.clk VPWR VGND sg13g2_buf_16
XFILLER_26_297 VPWR VGND sg13g2_fill_2
XFILLER_41_278 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3930_ heichips25_sap3/net435 VGND VPWR heichips25_sap3/_0071_ heichips25_sap3__3930_/Q
+ clkload23/A sg13g2_dfrbpq_1
XFILLER_10_643 VPWR VGND sg13g2_fill_1
XFILLER_5_102 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3861_ heichips25_sap3/net1019 VPWR heichips25_sap3/_1357_ VGND heichips25_sap3/net1064
+ heichips25_sap3/_1366_ sg13g2_o21ai_1
Xheichips25_sap3__2812_ VPWR VGND heichips25_sap3/_0456_ heichips25_sap3/net70 heichips25_sap3/_0455_
+ heichips25_sap3/_0212_ heichips25_sap3/_0457_ heichips25_sap3/net158 sg13g2_a221oi_1
Xheichips25_sap3__3792_ VPWR VGND heichips25_sap3/_1301_ heichips25_sap3/net339 heichips25_sap3/_1297_
+ heichips25_sap3/_1375_ heichips25_sap3/_1302_ heichips25_sap3/net290 sg13g2_a221oi_1
XFILLER_2_842 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2743_ heichips25_sap3/net288 heichips25_sap3__3915_/Q heichips25_sap3/_0389_
+ VPWR VGND sg13g2_nor2b_1
XFILLER_2_853 VPWR VGND sg13g2_decap_4
XFILLER_49_312 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2674_ heichips25_sap3/_1451_ heichips25_sap3/net237 heichips25_sap3/_1443_
+ heichips25_sap3/_0002_ VPWR VGND sg13g2_nand3_1
XFILLER_18_732 VPWR VGND sg13g2_fill_1
XFILLER_45_573 VPWR VGND sg13g2_decap_4
XFILLER_45_551 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3226_ heichips25_sap3/_0839_ heichips25_sap3__3965_/Q heichips25_sap3/net145
+ VPWR VGND sg13g2_nand2_1
XFILLER_27_90 VPWR VGND sg13g2_fill_1
XFILLER_17_275 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3157_ heichips25_sap3/_0666_ heichips25_sap3/_0679_ heichips25_sap3/_0697_
+ heichips25_sap3/_0770_ VPWR VGND sg13g2_nor3_1
Xheichips25_sap3__2108_ heichips25_sap3/net260 heichips25_sap3/net258 heichips25_sap3/_1529_
+ VPWR VGND heichips25_sap3/net272 sg13g2_nand3b_1
Xheichips25_sap3__3088_ heichips25_sap3/_0700_ VPWR heichips25_sap3/_0701_ VGND heichips25_sap3/net243
+ heichips25_sap3/_0307_ sg13g2_o21ai_1
XFILLER_20_429 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2039_ heichips25_sap3/_1460_ heichips25_sap3/net253 heichips25_sap3/net252
+ VPWR VGND sg13g2_nand2_1
XFILLER_9_496 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2714_ heichips25_can_lehmann_fsm/net485 VPWR heichips25_can_lehmann_fsm/_0823_
+ VGND heichips25_can_lehmann_fsm/net1039 heichips25_can_lehmann_fsm/net378 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2645_ VGND VPWR heichips25_can_lehmann_fsm/_0886_ heichips25_can_lehmann_fsm/net401
+ heichips25_can_lehmann_fsm/_0222_ heichips25_can_lehmann_fsm/_0788_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2576_ heichips25_can_lehmann_fsm/net482 VPWR heichips25_can_lehmann_fsm/_0754_
+ VGND heichips25_can_lehmann_fsm/net1038 heichips25_can_lehmann_fsm/net370 sg13g2_o21ai_1
XFILLER_23_15 VPWR VGND sg13g2_decap_4
XFILLER_23_267 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__3059_ net718 VGND VPWR heichips25_can_lehmann_fsm/net1133
+ heichips25_can_lehmann_fsm__3059_/Q clknet_leaf_14_clk sg13g2_dfrbpq_1
XFILLER_24_1025 VPWR VGND sg13g2_decap_4
XFILLER_47_838 VPWR VGND sg13g2_fill_2
XFILLER_46_315 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2390_ heichips25_sap3/_1809_ heichips25_sap3/net75 heichips25_sap3__3985_/Q
+ heichips25_sap3/net85 heichips25_sap3__3953_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_46_326 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__4060_ heichips25_sap3/net462 VGND VPWR heichips25_sap3/_0018_ heichips25_sap3/_0008_
+ clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_15_724 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3011_ heichips25_sap3/_0631_ VPWR heichips25_sap3/_0064_ VGND heichips25_sap3/net231
+ heichips25_sap3/_0212_ sg13g2_o21ai_1
XFILLER_15_768 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2823__561 VPWR VGND net560 sg13g2_tiehi
XFILLER_11_985 VPWR VGND sg13g2_fill_2
XFILLER_6_433 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3913_ heichips25_sap3/net454 VGND VPWR heichips25_sap3/_0054_ heichips25_sap3__3913_/Q
+ clkload25/A sg13g2_dfrbpq_1
Xheichips25_sap3__3844_ heichips25_sap3/net1223 VPWR heichips25_sap3/_1345_ VGND heichips25_sap3/_0018_
+ heichips25_sap3/_1260_ sg13g2_o21ai_1
XFILLER_6_477 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3775_ heichips25_sap3/_1286_ VPWR heichips25_sap3/_0173_ VGND heichips25_sap3/_1427_
+ heichips25_sap3__4062_/D sg13g2_o21ai_1
Xheichips25_sap3__2726_ heichips25_sap3__3915_/Q heichips25_sap3/net288 heichips25_sap3/_0372_
+ VPWR VGND sg13g2_xor2_1
Xheichips25_sap3__2657_ heichips25_sap3/_0324_ heichips25_sap3/_1679_ heichips25_sap3/_0323_
+ VPWR VGND sg13g2_nand2_1
XFILLER_49_142 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2588_ VGND VPWR heichips25_sap3/net156 heichips25_sap3/_0260_ heichips25_sap3/_0261_
+ heichips25_sap3/_0259_ sg13g2_a21oi_1
XFILLER_18_540 VPWR VGND sg13g2_fill_1
XFILLER_45_381 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3209_ heichips25_sap3/_0717_ heichips25_sap3/net151 heichips25_sap3__4019_/Q
+ heichips25_sap3/_0822_ VPWR VGND sg13g2_nand3_1
Xheichips25_can_lehmann_fsm__2430_ heichips25_can_lehmann_fsm/net481 VPWR heichips25_can_lehmann_fsm/_0681_
+ VGND heichips25_can_lehmann_fsm/net973 heichips25_can_lehmann_fsm/net412 sg13g2_o21ai_1
XFILLER_21_716 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2361_ VGND VPWR heichips25_can_lehmann_fsm/_0961_ heichips25_can_lehmann_fsm/net387
+ heichips25_can_lehmann_fsm/_0080_ heichips25_can_lehmann_fsm/_0646_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2292_ VGND VPWR heichips25_can_lehmann_fsm/_1051_ heichips25_can_lehmann_fsm/_0603_
+ heichips25_can_lehmann_fsm/_0604_ heichips25_can_lehmann_fsm/net171 sg13g2_a21oi_1
XFILLER_9_293 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm_fanout303 heichips25_can_lehmann_fsm/net304 heichips25_can_lehmann_fsm/net303
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout314 heichips25_can_lehmann_fsm/net316 heichips25_can_lehmann_fsm/net314
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout325 heichips25_can_lehmann_fsm/net326 heichips25_can_lehmann_fsm/net325
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout347 heichips25_can_lehmann_fsm/net1269 heichips25_can_lehmann_fsm/net347
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout336 heichips25_can_lehmann_fsm/_1001_ heichips25_can_lehmann_fsm/net336
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm__2991__661 VPWR VGND net660 sg13g2_tiehi
Xheichips25_can_lehmann_fsm_fanout369 heichips25_can_lehmann_fsm/net371 heichips25_can_lehmann_fsm/net369
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout358 heichips25_can_lehmann_fsm/net361 heichips25_can_lehmann_fsm/net358
+ VPWR VGND sg13g2_buf_1
XFILLER_18_48 VPWR VGND sg13g2_fill_1
XFILLER_34_36 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2628_ heichips25_can_lehmann_fsm/net477 VPWR heichips25_can_lehmann_fsm/_0780_
+ VGND heichips25_can_lehmann_fsm/net963 heichips25_can_lehmann_fsm/net368 sg13g2_o21ai_1
XFILLER_11_215 VPWR VGND sg13g2_fill_1
XFILLER_11_237 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2559_ VGND VPWR heichips25_can_lehmann_fsm/_0908_ heichips25_can_lehmann_fsm/net430
+ heichips25_can_lehmann_fsm/_0179_ heichips25_can_lehmann_fsm/_0745_ sg13g2_a21oi_1
Xclkload2 clknet_leaf_13_clk clkload2/X VPWR VGND sg13g2_buf_8
XFILLER_4_959 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3560_ heichips25_sap3__3962_/Q heichips25_sap3/_1083_ heichips25_sap3/net56
+ heichips25_sap3/_0103_ VPWR VGND sg13g2_mux2_1
Xheichips25_can_lehmann_fsm__2970__745 VPWR VGND net744 sg13g2_tiehi
Xheichips25_sap3__2511_ heichips25_sap3__3898_/Q heichips25_sap3/net215 heichips25_sap3/_1923_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__3491_ heichips25_sap3/_1088_ heichips25_sap3/net108 heichips25_sap3/net131
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__2442_ heichips25_sap3/_1857_ heichips25_sap3/net75 heichips25_sap3__3991_/Q
+ heichips25_sap3/net90 heichips25_sap3__3943_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_19_337 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2373_ heichips25_sap3/_1794_ heichips25_sap3/net75 heichips25_sap3__3994_/Q
+ heichips25_sap3/net81 heichips25_sap3__3978_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_28_871 VPWR VGND sg13g2_fill_2
XFILLER_28_893 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__4043_ heichips25_sap3/net460 VGND VPWR heichips25_sap3/_0184_ heichips25_sap3__4043_/Q
+ clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_15_576 VPWR VGND sg13g2_decap_8
XFILLER_30_546 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_hold970 heichips25_can_lehmann_fsm__2944_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net969 sg13g2_dlygate4sd3_1
XFILLER_24_80 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm_hold981 heichips25_can_lehmann_fsm__2860_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net980 sg13g2_dlygate4sd3_1
XFILLER_7_731 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm_hold992 heichips25_can_lehmann_fsm/_0244_ VPWR VGND heichips25_can_lehmann_fsm/net991
+ sg13g2_dlygate4sd3_1
XFILLER_6_274 VPWR VGND sg13g2_decap_8
Xclkbuf_5_24__f_heichips25_sap3\_sap_3_inst.alu_inst.clk heichips25_sap3__4005_/CLK
+ clknet_4_12_0_heichips25_sap3\/sap_3_inst.alu_inst.clk VPWR VGND sg13g2_buf_16
Xheichips25_sap3__3827_ VPWR VGND heichips25_sap3__3953_/Q heichips25_sap3/_1332_
+ heichips25_sap3/_1282_ heichips25_sap3__4009_/Q heichips25_sap3/_1333_ heichips25_sap3/_1278_
+ sg13g2_a221oi_1
Xheichips25_sap3__3758_ heichips25_sap3/_1260_ heichips25_sap3/_1264_ heichips25_sap3/_1270_
+ VPWR VGND sg13g2_nor2_1
XFILLER_3_970 VPWR VGND sg13g2_decap_8
XFILLER_34_4 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2709_ heichips25_sap3/_0355_ heichips25_sap3/net280 heichips25_sap3__3919_/Q
+ VPWR VGND sg13g2_xnor2_1
Xheichips25_sap3__3689_ heichips25_sap3/net111 heichips25_sap3/_0984_ heichips25_sap3/_1069_
+ heichips25_sap3/_1137_ heichips25_sap3/_1226_ VPWR VGND sg13g2_nor4_1
Xheichips25_can_lehmann_fsm__1930_ heichips25_can_lehmann_fsm/_0293_ heichips25_can_lehmann_fsm/_1162_
+ heichips25_can_lehmann_fsm/_0292_ VPWR VGND sg13g2_nand2b_1
Xheichips25_can_lehmann_fsm__1861_ heichips25_can_lehmann_fsm/_1174_ heichips25_can_lehmann_fsm/_0984_
+ heichips25_can_lehmann_fsm/_1165_ heichips25_can_lehmann_fsm/_1177_ VPWR VGND sg13g2_mux2_1
X_26_ net511 uio_oe_sap3\[4\] net506 net23 VPWR VGND sg13g2_mux2_1
Xheichips25_can_lehmann_fsm__1792_ heichips25_can_lehmann_fsm/_1108_ heichips25_can_lehmann_fsm/_1107_
+ heichips25_can_lehmann_fsm/_1104_ VPWR VGND sg13g2_nand2b_1
Xheichips25_sap3_fanout218 heichips25_sap3/_1724_ heichips25_sap3/net218 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout229 heichips25_sap3/_1497_ heichips25_sap3/net229 VPWR VGND
+ sg13g2_buf_1
Xheichips25_can_lehmann_fsm__2413_ VGND VPWR heichips25_can_lehmann_fsm/_0946_ heichips25_can_lehmann_fsm/net380
+ heichips25_can_lehmann_fsm/_0106_ heichips25_can_lehmann_fsm/_0672_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2344_ heichips25_can_lehmann_fsm/net494 VPWR heichips25_can_lehmann_fsm/_0638_
+ VGND heichips25_can_lehmann_fsm/net1034 heichips25_can_lehmann_fsm/net367 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2275_ VGND VPWR heichips25_can_lehmann_fsm/net207 heichips25_can_lehmann_fsm/_0589_
+ heichips25_can_lehmann_fsm/_0050_ heichips25_can_lehmann_fsm/_0590_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm_fanout199 heichips25_can_lehmann_fsm/net200 heichips25_can_lehmann_fsm/net199
+ VPWR VGND sg13g2_buf_1
XFILLER_0_417 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_fanout188 heichips25_can_lehmann_fsm/net190 heichips25_can_lehmann_fsm/net188
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout177 heichips25_can_lehmann_fsm/net180 heichips25_can_lehmann_fsm/net177
+ VPWR VGND sg13g2_buf_1
XFILLER_28_101 VPWR VGND sg13g2_decap_8
XFILLER_21_1028 VPWR VGND sg13g2_fill_1
XFILLER_45_57 VPWR VGND sg13g2_fill_1
XFILLER_40_822 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2991_ heichips25_sap3/_0621_ heichips25_sap3__3914_/Q heichips25_sap3/_0607_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__1942_ VPWR heichips25_sap3/_1368_ heichips25_sap3__3934_/Q VGND
+ sg13g2_inv_1
XFILLER_3_233 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3612_ heichips25_sap3/_1178_ heichips25_sap3__3978_/Q heichips25_sap3/_1171_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__3543_ heichips25_sap3/net107 heichips25_sap3/_1131_ heichips25_sap3/_1132_
+ heichips25_sap3/_1133_ VPWR VGND sg13g2_nor3_1
Xheichips25_sap3__3474_ heichips25_sap3/_0863_ heichips25_sap3/_0995_ heichips25_sap3/_1074_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__2425_ heichips25_sap3/_1842_ heichips25_sap3/net84 heichips25_sap3__3968_/Q
+ heichips25_sap3/net91 heichips25_sap3__3944_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_47_498 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2356_ heichips25_sap3/net256 heichips25_sap3/_1480_ heichips25_sap3/_1492_
+ heichips25_sap3/_1777_ VPWR VGND sg13g2_nor3_1
XFILLER_19_189 VPWR VGND sg13g2_fill_1
XFILLER_34_137 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2287_ VGND VPWR heichips25_sap3/net270 heichips25_sap3/_1649_ heichips25_sap3/_1708_
+ heichips25_sap3/_1453_ sg13g2_a21oi_1
Xheichips25_sap3__4026_ heichips25_sap3/net445 VGND VPWR heichips25_sap3/_0167_ heichips25_sap3__4026_/Q
+ clkload22/A sg13g2_dfrbpq_1
XFILLER_30_387 VPWR VGND sg13g2_fill_2
XFILLER_7_550 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2060_ heichips25_can_lehmann_fsm/net1255 heichips25_can_lehmann_fsm/net182
+ heichips25_can_lehmann_fsm/_0408_ VPWR VGND sg13g2_nor2_1
XFILLER_39_911 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2962_ net776 VGND VPWR heichips25_can_lehmann_fsm/_0187_
+ heichips25_can_lehmann_fsm__2962_/Q clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_39_977 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2893_ net709 VGND VPWR heichips25_can_lehmann_fsm/_0118_
+ heichips25_can_lehmann_fsm__2893_/Q clknet_leaf_18_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1913_ heichips25_can_lehmann_fsm/_1226_ heichips25_can_lehmann_fsm/_0895_
+ heichips25_can_lehmann_fsm/net349 VPWR VGND sg13g2_nand2_1
Xheichips25_can_lehmann_fsm__1844_ heichips25_can_lehmann_fsm/_1141_ heichips25_can_lehmann_fsm/_1108_
+ heichips25_can_lehmann_fsm/_1158_ heichips25_can_lehmann_fsm/_1160_ VPWR VGND sg13g2_a21o_1
XFILLER_26_616 VPWR VGND sg13g2_fill_1
X_09_ uo_out_fsm\[3\] uo_out_sap3\[3\] net507 net38 VPWR VGND sg13g2_mux2_1
XFILLER_41_619 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm_hold1105 heichips25_can_lehmann_fsm/_0179_ VPWR VGND heichips25_can_lehmann_fsm/net1104
+ sg13g2_dlygate4sd3_1
XFILLER_34_671 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1775_ heichips25_can_lehmann_fsm/_1091_ heichips25_can_lehmann_fsm/net332
+ heichips25_can_lehmann_fsm__3037_/Q heichips25_can_lehmann_fsm/net317 heichips25_can_lehmann_fsm__2989_/Q
+ VPWR VGND sg13g2_a22oi_1
XFILLER_22_800 VPWR VGND sg13g2_fill_1
XFILLER_40_129 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_hold1116 heichips25_can_lehmann_fsm__2848_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1115 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1138 heichips25_can_lehmann_fsm__3060_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1137 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1127 heichips25_can_lehmann_fsm__2877_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1126 sg13g2_dlygate4sd3_1
Xheichips25_sap3_hold836 heichips25_sap3__4031_/Q VPWR VGND heichips25_sap3/net835
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1149 heichips25_can_lehmann_fsm__3058_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1148 sg13g2_dlygate4sd3_1
XFILLER_5_509 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2327_ VGND VPWR heichips25_can_lehmann_fsm/_0970_ heichips25_can_lehmann_fsm/net403
+ heichips25_can_lehmann_fsm/_0063_ heichips25_can_lehmann_fsm/_0629_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2258_ heichips25_can_lehmann_fsm/net327 VPWR heichips25_can_lehmann_fsm/_0577_
+ VGND heichips25_can_lehmann_fsm__2822_/Q heichips25_can_lehmann_fsm/net206 sg13g2_o21ai_1
Xheichips25_sap3_fanout57 heichips25_sap3/net58 heichips25_sap3/net57 VPWR VGND sg13g2_buf_1
Xheichips25_sap3_fanout68 heichips25_sap3/_0883_ heichips25_sap3/net68 VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm__2189_ heichips25_can_lehmann_fsm/net325 VPWR heichips25_can_lehmann_fsm/_0523_
+ VGND heichips25_can_lehmann_fsm/net1210 heichips25_can_lehmann_fsm/net160 sg13g2_o21ai_1
Xoutput37 net37 uo_out[2] VPWR VGND sg13g2_buf_1
Xheichips25_sap3_fanout79 heichips25_sap3/_1741_ heichips25_sap3/net79 VPWR VGND sg13g2_buf_1
Xoutput26 net26 uio_oe[7] VPWR VGND sg13g2_buf_1
Xheichips25_sap3__2210_ heichips25_sap3/_1482_ heichips25_sap3/net223 heichips25_sap3/_1631_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__3190_ heichips25_sap3/_0803_ heichips25_sap3/net139 heichips25_sap3__3983_/Q
+ heichips25_sap3/net142 heichips25_sap3__3991_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2141_ VGND VPWR heichips25_sap3/_1544_ heichips25_sap3/_1561_ heichips25_sap3/_1562_
+ heichips25_sap3/_1558_ sg13g2_a21oi_1
XFILLER_25_660 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2072_ heichips25_sap3/_1493_ heichips25_sap3/_1485_ heichips25_sap3/_1491_
+ VPWR VGND sg13g2_nand2_1
XFILLER_12_310 VPWR VGND sg13g2_decap_8
XFILLER_8_325 VPWR VGND sg13g2_fill_1
XFILLER_8_358 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2974_ heichips25_sap3/_0610_ heichips25_sap3__3908_/Q heichips25_sap3/_0607_
+ VPWR VGND sg13g2_nand2_1
XFILLER_21_70 VPWR VGND sg13g2_fill_1
XFILLER_4_553 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3526_ heichips25_sap3/net120 VPWR heichips25_sap3/_1118_ VGND heichips25_sap3/net828
+ heichips25_sap3/_1088_ sg13g2_o21ai_1
XFILLER_11_6 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3457_ heichips25_sap3/_0903_ heichips25_sap3/net122 uio_out_sap3\[1\]
+ heichips25_sap3/_1061_ VPWR VGND sg13g2_a21o_1
XFILLER_47_251 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2408_ heichips25_sap3/_1825_ heichips25_sap3/net84 heichips25_sap3__3960_/Q
+ heichips25_sap3/net87 heichips25_sap3__3944_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3388_ VGND VPWR heichips25_sap3/net123 heichips25_sap3/_0995_ heichips25_sap3/_0996_
+ heichips25_sap3/_0863_ sg13g2_a21oi_1
XFILLER_35_435 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2339_ VGND VPWR heichips25_sap3/net227 heichips25_sap3/_1623_ heichips25_sap3/_1760_
+ heichips25_sap3/net223 sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__1560_ VPWR heichips25_can_lehmann_fsm/_0884_ heichips25_can_lehmann_fsm/net860
+ VGND sg13g2_inv_1
Xheichips25_sap3__4009_ heichips25_sap3/net444 VGND VPWR heichips25_sap3/_0150_ heichips25_sap3__4009_/Q
+ heichips25_sap3__4009_/CLK sg13g2_dfrbpq_1
XFILLER_31_652 VPWR VGND sg13g2_decap_8
XFILLER_31_696 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2112_ heichips25_can_lehmann_fsm/_0449_ heichips25_can_lehmann_fsm/_0450_
+ heichips25_can_lehmann_fsm/_0448_ heichips25_can_lehmann_fsm/_0451_ VPWR VGND sg13g2_nand3_1
Xheichips25_can_lehmann_fsm__2043_ net11 heichips25_can_lehmann_fsm/_1215_ heichips25_can_lehmann_fsm/_0392_
+ VPWR VGND sg13g2_and2_1
Xheichips25_can_lehmann_fsm__2945_ net555 VGND VPWR heichips25_can_lehmann_fsm/_0170_
+ heichips25_can_lehmann_fsm__2945_/Q clknet_leaf_21_clk sg13g2_dfrbpq_1
XFILLER_26_15 VPWR VGND sg13g2_decap_8
XFILLER_26_26 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2876_ net743 VGND VPWR heichips25_can_lehmann_fsm/net1111
+ heichips25_can_lehmann_fsm__2876_/Q clknet_leaf_1_clk sg13g2_dfrbpq_1
XFILLER_42_939 VPWR VGND sg13g2_fill_2
XFILLER_42_928 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1827_ heichips25_can_lehmann_fsm__3045_/Q heichips25_can_lehmann_fsm/net343
+ heichips25_can_lehmann_fsm/_1143_ VPWR VGND sg13g2_nor2b_1
XFILLER_26_468 VPWR VGND sg13g2_fill_2
XFILLER_41_449 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1758_ uo_out_fsm\[4\] heichips25_can_lehmann_fsm/_1076_
+ heichips25_can_lehmann_fsm/_1077_ VPWR VGND sg13g2_nand2_1
XFILLER_10_803 VPWR VGND sg13g2_fill_1
XFILLER_10_836 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__1689_ heichips25_can_lehmann_fsm/_1013_ heichips25_can_lehmann_fsm/net294
+ heichips25_can_lehmann_fsm__2970_/Q heichips25_can_lehmann_fsm/net310 heichips25_can_lehmann_fsm__3018_/Q
+ VPWR VGND sg13g2_a22oi_1
XFILLER_10_847 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2690_ heichips25_sap3/_0336_ heichips25_sap3__3898_/Q heichips25_sap3/_0335_
+ VPWR VGND sg13g2_nand2b_1
XFILLER_49_505 VPWR VGND sg13g2_decap_8
XFILLER_18_903 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3311_ VGND VPWR heichips25_sap3/_1375_ heichips25_sap3/net127 heichips25_sap3/_0922_
+ heichips25_sap3/_0921_ sg13g2_a21oi_1
XFILLER_18_925 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3242_ heichips25_sap3/net61 heichips25_sap3/_0841_ heichips25_sap3/_0819_
+ heichips25_sap3/_0855_ VPWR VGND heichips25_sap3/_0852_ sg13g2_nand4_1
Xheichips25_sap3__3173_ heichips25_sap3/_0782_ heichips25_sap3/_0785_ heichips25_sap3/_0786_
+ VPWR VGND sg13g2_nor2_1
XFILLER_17_468 VPWR VGND sg13g2_fill_2
XFILLER_33_906 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2124_ heichips25_sap3/_1545_ heichips25_sap3/net229 heichips25_sap3/_1544_
+ VPWR VGND sg13g2_nand2_1
XFILLER_16_81 VPWR VGND sg13g2_fill_1
XFILLER_40_471 VPWR VGND sg13g2_fill_2
XFILLER_40_460 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2055_ heichips25_sap3/_1444_ heichips25_sap3/_1475_ heichips25_sap3/_1476_
+ VPWR VGND sg13g2_nor2_1
XFILLER_12_162 VPWR VGND sg13g2_decap_8
XFILLER_5_840 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2957_ VPWR VGND heichips25_sap3/_0381_ heichips25_sap3/_0594_ heichips25_sap3/_0445_
+ heichips25_sap3/net276 heichips25_sap3/_0595_ heichips25_sap3/_0417_ sg13g2_a221oi_1
Xheichips25_sap3__2888_ heichips25_sap3/net64 heichips25_sap3/_0528_ heichips25_sap3/_0529_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_can_lehmann_fsm__2833__541 VPWR VGND net540 sg13g2_tiehi
XFILLER_48_571 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3509_ VGND VPWR heichips25_sap3/_1104_ heichips25_sap3/_0914_ heichips25_sap3/net119
+ sg13g2_or2_1
Xheichips25_can_lehmann_fsm__2730_ heichips25_can_lehmann_fsm/net466 VPWR heichips25_can_lehmann_fsm/_0831_
+ VGND heichips25_can_lehmann_fsm__3039_/Q heichips25_can_lehmann_fsm/net356 sg13g2_o21ai_1
XFILLER_35_265 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2661_ VGND VPWR heichips25_can_lehmann_fsm/_0880_ heichips25_can_lehmann_fsm/net384
+ heichips25_can_lehmann_fsm/_0230_ heichips25_can_lehmann_fsm/_0796_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__1612_ VPWR heichips25_can_lehmann_fsm/_0936_ heichips25_can_lehmann_fsm/net913
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__2909__678 VPWR VGND net677 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2592_ heichips25_can_lehmann_fsm/net468 VPWR heichips25_can_lehmann_fsm/_0762_
+ VGND heichips25_can_lehmann_fsm__2970_/Q heichips25_can_lehmann_fsm/net360 sg13g2_o21ai_1
Xclkbuf_leaf_15_clk clknet_2_2__leaf_clk clknet_leaf_15_clk VPWR VGND sg13g2_buf_8
Xheichips25_can_lehmann_fsm__1543_ VPWR heichips25_can_lehmann_fsm/_0867_ heichips25_can_lehmann_fsm/net951
+ VGND sg13g2_inv_1
XFILLER_32_983 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__3055__671 VPWR VGND net670 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2026_ heichips25_can_lehmann_fsm/net321 VPWR heichips25_can_lehmann_fsm/_0378_
+ VGND heichips25_can_lehmann_fsm/net1246 heichips25_can_lehmann_fsm/net178 sg13g2_o21ai_1
XFILLER_39_560 VPWR VGND sg13g2_fill_1
XFILLER_2_1014 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2928_ net623 VGND VPWR heichips25_can_lehmann_fsm/net1063
+ heichips25_can_lehmann_fsm__2928_/Q clknet_leaf_13_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2859_ net777 VGND VPWR heichips25_can_lehmann_fsm/net943
+ heichips25_can_lehmann_fsm__2859_/Q clknet_leaf_10_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2966__761 VPWR VGND net760 sg13g2_tiehi
XFILLER_6_637 VPWR VGND sg13g2_fill_2
XFILLER_5_136 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3860_ VGND VPWR heichips25_sap3/net1065 heichips25_sap3/_1346_ heichips25_sap3/_0188_
+ heichips25_sap3/net1072 sg13g2_a21oi_1
Xheichips25_sap3__2811_ VGND VPWR heichips25_sap3__3907_/Q heichips25_sap3/net204
+ heichips25_sap3/_0456_ heichips25_sap3/net158 sg13g2_a21oi_1
Xheichips25_sap3__3791_ VPWR VGND heichips25_sap3__4021_/Q heichips25_sap3/_1300_
+ heichips25_sap3/_1270_ heichips25_sap3__3997_/Q heichips25_sap3/_1301_ heichips25_sap3/_1265_
+ sg13g2_a221oi_1
XFILLER_2_810 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2742_ heichips25_sap3/net283 heichips25_sap3__3918_/Q heichips25_sap3/_0388_
+ VPWR VGND sg13g2_nor2b_1
Xheichips25_sap3__2673_ VPWR VGND heichips25_sap3/_1751_ heichips25_sap3/_1593_ heichips25_sap3/_1747_
+ heichips25_sap3/_1420_ uio_oe_sap3\[7\] heichips25_sap3/net91 sg13g2_a221oi_1
XFILLER_49_324 VPWR VGND sg13g2_decap_8
XFILLER_49_368 VPWR VGND sg13g2_decap_8
XFILLER_17_210 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3225_ heichips25_sap3/_0680_ heichips25_sap3/net152 heichips25_sap3__3941_/Q
+ heichips25_sap3/_0838_ VPWR VGND sg13g2_nand3_1
XFILLER_18_799 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3156_ heichips25_sap3/_0769_ heichips25_sap3/net138 heichips25_sap3__3971_/Q
+ heichips25_sap3/net140 heichips25_sap3__3979_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3087_ heichips25_sap3/_1468_ heichips25_sap3/_1552_ heichips25_sap3/_0700_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__2107_ heichips25_sap3/_1503_ heichips25_sap3/_1522_ heichips25_sap3/_1526_
+ heichips25_sap3/_1528_ VPWR VGND sg13g2_nor3_1
XFILLER_13_482 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2038_ heichips25_sap3/net253 heichips25_sap3/net252 heichips25_sap3/_1459_
+ VPWR VGND sg13g2_and2_1
Xheichips25_sap3__3989_ heichips25_sap3/net456 VGND VPWR heichips25_sap3/_0130_ heichips25_sap3__3989_/Q
+ heichips25_sap3__4003_/CLK sg13g2_dfrbpq_1
Xclkbuf_leaf_4_clk clknet_2_1__leaf_clk clknet_leaf_4_clk VPWR VGND sg13g2_buf_8
XFILLER_48_390 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2713_ VGND VPWR heichips25_can_lehmann_fsm/_0867_ heichips25_can_lehmann_fsm/net417
+ heichips25_can_lehmann_fsm/_0256_ heichips25_can_lehmann_fsm/_0822_ sg13g2_a21oi_1
XFILLER_17_1000 VPWR VGND sg13g2_fill_2
XFILLER_23_235 VPWR VGND sg13g2_fill_1
XFILLER_24_769 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2644_ heichips25_can_lehmann_fsm/net473 VPWR heichips25_can_lehmann_fsm/_0788_
+ VGND heichips25_can_lehmann_fsm/net855 heichips25_can_lehmann_fsm/net401 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2575_ VGND VPWR heichips25_can_lehmann_fsm/_0904_ heichips25_can_lehmann_fsm/net409
+ heichips25_can_lehmann_fsm/_0187_ heichips25_can_lehmann_fsm/_0753_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__3018__739 VPWR VGND net738 sg13g2_tiehi
XFILLER_2_117 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__3058_ net782 VGND VPWR heichips25_can_lehmann_fsm/_0283_
+ heichips25_can_lehmann_fsm__3058_/Q clknet_leaf_16_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2009_ heichips25_can_lehmann_fsm/_0363_ heichips25_can_lehmann_fsm/_1070_
+ heichips25_can_lehmann_fsm/_0362_ VPWR VGND sg13g2_nand2_1
XFILLER_48_35 VPWR VGND sg13g2_fill_2
XFILLER_46_338 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3010_ heichips25_sap3/_0631_ heichips25_sap3/net273 heichips25_sap3/net231
+ VPWR VGND sg13g2_nand2_1
XFILLER_14_213 VPWR VGND sg13g2_fill_1
XFILLER_42_588 VPWR VGND sg13g2_fill_1
XFILLER_42_577 VPWR VGND sg13g2_fill_2
XFILLER_23_791 VPWR VGND sg13g2_decap_8
XFILLER_11_953 VPWR VGND sg13g2_decap_8
XFILLER_11_964 VPWR VGND sg13g2_fill_1
XFILLER_6_445 VPWR VGND sg13g2_fill_1
XFILLER_6_412 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3912_ heichips25_sap3/net454 VGND VPWR heichips25_sap3/_0053_ heichips25_sap3__3912_/Q
+ clkload25/A sg13g2_dfrbpq_1
XFILLER_13_82 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3843_ heichips25_sap3/_1344_ VPWR heichips25_sap3/_0183_ VGND heichips25_sap3/_0018_
+ heichips25_sap3/_1267_ sg13g2_o21ai_1
XFILLER_6_456 VPWR VGND sg13g2_decap_8
XFILLER_6_489 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3774_ heichips25_sap3/_1285_ VPWR heichips25_sap3/_1286_ VGND heichips25_sap3/_1269_
+ heichips25_sap3/_1284_ sg13g2_o21ai_1
Xheichips25_sap3__2725_ heichips25_sap3/_0348_ VPWR heichips25_sap3/_0371_ VGND heichips25_sap3/_0347_
+ heichips25_sap3/_0370_ sg13g2_o21ai_1
Xheichips25_sap3__2656_ heichips25_sap3/_0323_ heichips25_sap3/_0321_ heichips25_sap3/_0322_
+ heichips25_sap3/net248 heichips25_sap3/_1447_ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2587_ heichips25_sap3/_0260_ heichips25_sap3__3890_/Q heichips25_sap3/_1788_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__3208_ heichips25_sap3/_0821_ heichips25_sap3__4003_/Q heichips25_sap3/net147
+ VPWR VGND sg13g2_nand2_1
XFILLER_33_555 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3139_ heichips25_sap3/_0717_ heichips25_sap3/net151 heichips25_sap3/_0752_
+ VPWR VGND sg13g2_and2_1
Xheichips25_can_lehmann_fsm__2360_ heichips25_can_lehmann_fsm/net500 VPWR heichips25_can_lehmann_fsm/_0646_
+ VGND heichips25_can_lehmann_fsm__2854_/Q heichips25_can_lehmann_fsm/net387 sg13g2_o21ai_1
XFILLER_20_216 VPWR VGND sg13g2_fill_1
XFILLER_9_261 VPWR VGND sg13g2_decap_8
Xclkload20 VPWR clkload20/Y clkload20/A VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__2291_ heichips25_can_lehmann_fsm/net1165 VPWR heichips25_can_lehmann_fsm/_0603_
+ VGND heichips25_can_lehmann_fsm__2828_/Q heichips25_can_lehmann_fsm/_1049_ sg13g2_o21ai_1
XFILLER_9_272 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_fanout304 heichips25_can_lehmann_fsm/_1000_ heichips25_can_lehmann_fsm/net304
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout326 heichips25_can_lehmann_fsm/net330 heichips25_can_lehmann_fsm/net326
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout337 heichips25_can_lehmann_fsm/_0998_ heichips25_can_lehmann_fsm/net337
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout348 heichips25_can_lehmann_fsm__2777_/Q heichips25_can_lehmann_fsm/net348
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout315 heichips25_can_lehmann_fsm/net316 heichips25_can_lehmann_fsm/net315
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout359 heichips25_can_lehmann_fsm/net360 heichips25_can_lehmann_fsm/net359
+ VPWR VGND sg13g2_buf_1
XFILLER_43_308 VPWR VGND sg13g2_decap_8
XFILLER_36_371 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2627_ VGND VPWR heichips25_can_lehmann_fsm/_0891_ heichips25_can_lehmann_fsm/net409
+ heichips25_can_lehmann_fsm/_0213_ heichips25_can_lehmann_fsm/_0779_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2558_ heichips25_can_lehmann_fsm/net500 VPWR heichips25_can_lehmann_fsm/_0745_
+ VGND heichips25_can_lehmann_fsm__2954_/Q heichips25_can_lehmann_fsm/net430 sg13g2_o21ai_1
XFILLER_11_249 VPWR VGND sg13g2_fill_1
Xclkload3 clkload3/Y clknet_leaf_21_clk VPWR VGND sg13g2_inv_2
Xheichips25_can_lehmann_fsm__2489_ VGND VPWR heichips25_can_lehmann_fsm/_0925_ heichips25_can_lehmann_fsm/net357
+ heichips25_can_lehmann_fsm/_0144_ heichips25_can_lehmann_fsm/_0710_ sg13g2_a21oi_1
XFILLER_3_404 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2510_ VPWR heichips25_sap3/_1922_ uio_out_sap3\[1\] VGND sg13g2_inv_1
Xheichips25_sap3__3490_ heichips25_sap3/net106 heichips25_sap3/_0882_ heichips25_sap3/_1087_
+ VPWR VGND sg13g2_nor2_1
Xclkbuf_5_7__f_heichips25_sap3\_sap_3_inst.alu_inst.clk clkload19/A clknet_4_3_0_heichips25_sap3\/sap_3_inst.alu_inst.clk
+ VPWR VGND sg13g2_buf_16
Xheichips25_sap3__2441_ heichips25_sap3/_1856_ heichips25_sap3/_1853_ heichips25_sap3/_1855_
+ heichips25_sap3/_1770_ net7 VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2372_ heichips25_sap3/_1793_ heichips25_sap3/net72 heichips25_sap3__3986_/Q
+ heichips25_sap3/net85 heichips25_sap3__3962_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_19_349 VPWR VGND sg13g2_decap_8
XFILLER_34_308 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__4042_ heichips25_sap3/net460 VGND VPWR heichips25_sap3/_0183_ heichips25_sap3__4042_/Q
+ clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_42_363 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm_hold971 heichips25_can_lehmann_fsm__2941_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net970 sg13g2_dlygate4sd3_1
XFILLER_24_70 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm_hold960 heichips25_can_lehmann_fsm__2974_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net959 sg13g2_dlygate4sd3_1
XFILLER_7_743 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm_hold982 heichips25_can_lehmann_fsm__2919_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net981 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold993 heichips25_can_lehmann_fsm__2931_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net992 sg13g2_dlygate4sd3_1
Xheichips25_sap3__3826_ heichips25_sap3/_1329_ heichips25_sap3/_1330_ heichips25_sap3/_1327_
+ heichips25_sap3/_1332_ VPWR VGND heichips25_sap3/_1331_ sg13g2_nand4_1
Xheichips25_sap3__3757_ heichips25_sap3/_1269_ heichips25_sap3/_1263_ heichips25_sap3/_1268_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__2708_ heichips25_sap3/net280 heichips25_sap3__3919_/Q heichips25_sap3/_0354_
+ VPWR VGND sg13g2_and2_1
XFILLER_27_4 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3688_ heichips25_sap3/_1225_ VPWR heichips25_sap3/_0147_ VGND heichips25_sap3/net112
+ heichips25_sap3/_1191_ sg13g2_o21ai_1
Xheichips25_sap3__2639_ VGND VPWR heichips25_sap3/net235 heichips25_sap3/_1569_ heichips25_sap3/_0306_
+ heichips25_sap3/_1565_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__1860_ heichips25_can_lehmann_fsm/_1176_ heichips25_can_lehmann_fsm/net471
+ net9 VPWR VGND sg13g2_nand2b_1
X_25_ net510 uio_oe_sap3\[3\] net506 net22 VPWR VGND sg13g2_mux2_1
Xheichips25_can_lehmann_fsm__1791_ heichips25_can_lehmann_fsm__2817_/Q heichips25_can_lehmann_fsm__2816_/Q
+ heichips25_can_lehmann_fsm__2815_/Q heichips25_can_lehmann_fsm__2814_/Q heichips25_can_lehmann_fsm/_1107_
+ VPWR VGND sg13g2_nor4_1
XFILLER_45_190 VPWR VGND sg13g2_decap_8
XFILLER_34_853 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2412_ heichips25_can_lehmann_fsm/net492 VPWR heichips25_can_lehmann_fsm/_0672_
+ VGND heichips25_can_lehmann_fsm__2880_/Q heichips25_can_lehmann_fsm/net380 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2343_ VGND VPWR heichips25_can_lehmann_fsm/_0966_ heichips25_can_lehmann_fsm/net406
+ heichips25_can_lehmann_fsm/_0071_ heichips25_can_lehmann_fsm/_0637_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2274_ heichips25_can_lehmann_fsm/net327 VPWR heichips25_can_lehmann_fsm/_0590_
+ VGND heichips25_can_lehmann_fsm/net1182 heichips25_can_lehmann_fsm/net207 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__3054__703 VPWR VGND net702 sg13g2_tiehi
XFILLER_20_28 VPWR VGND sg13g2_decap_8
XFILLER_1_919 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm_fanout178 heichips25_can_lehmann_fsm/net180 heichips25_can_lehmann_fsm/net178
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout189 heichips25_can_lehmann_fsm/net190 heichips25_can_lehmann_fsm/net189
+ VPWR VGND sg13g2_buf_1
XFILLER_44_606 VPWR VGND sg13g2_fill_1
XFILLER_28_157 VPWR VGND sg13g2_decap_8
XFILLER_25_820 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1989_ VGND VPWR heichips25_can_lehmann_fsm__2785_/Q heichips25_can_lehmann_fsm/net189
+ heichips25_can_lehmann_fsm/_0346_ heichips25_can_lehmann_fsm/net194 sg13g2_a21oi_1
XFILLER_43_138 VPWR VGND sg13g2_fill_1
XFILLER_25_853 VPWR VGND sg13g2_fill_2
XFILLER_24_363 VPWR VGND sg13g2_decap_8
XFILLER_25_864 VPWR VGND sg13g2_fill_2
XFILLER_40_834 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2990_ heichips25_sap3/_0054_ heichips25_sap3/_0619_ heichips25_sap3/_0620_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__1941_ VPWR heichips25_sap3/_1367_ heichips25_sap3/net282 VGND sg13g2_inv_1
XFILLER_3_245 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3611_ heichips25_sap3/_1083_ heichips25_sap3/_1128_ heichips25_sap3/_1177_
+ VPWR VGND sg13g2_nor2_1
XFILLER_3_256 VPWR VGND sg13g2_fill_1
XFILLER_10_50 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3542_ net47 uio_oe_sap3\[7\] heichips25_sap3/_1087_ heichips25_sap3/_1132_
+ VPWR VGND sg13g2_mux2_1
XFILLER_47_411 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3473_ heichips25_sap3/_1003_ heichips25_sap3/net121 uio_out_sap3\[5\]
+ heichips25_sap3/_1073_ VPWR VGND sg13g2_a21o_1
XFILLER_0_985 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2424_ heichips25_sap3/_1841_ heichips25_sap3/_1740_ heichips25_sap3__3976_/Q
+ heichips25_sap3/net88 heichips25_sap3__3952_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_19_70 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2355_ VGND VPWR heichips25_sap3/_1517_ heichips25_sap3/_1549_ heichips25_sap3/_1776_
+ heichips25_sap3/net223 sg13g2_a21oi_1
XFILLER_16_842 VPWR VGND sg13g2_decap_8
XFILLER_43_661 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2286_ heichips25_sap3/_1706_ heichips25_sap3/_1641_ heichips25_sap3/_1707_
+ VPWR VGND heichips25_sap3/_1705_ sg13g2_nand3b_1
XFILLER_15_330 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__4025_ heichips25_sap3/net459 VGND VPWR heichips25_sap3/_0166_ heichips25_sap3__4025_/Q
+ clkload29/A sg13g2_dfrbpq_1
XFILLER_35_80 VPWR VGND sg13g2_fill_2
XFILLER_31_823 VPWR VGND sg13g2_fill_2
XFILLER_31_834 VPWR VGND sg13g2_decap_4
XFILLER_30_355 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3809_ VPWR VGND heichips25_sap3__3999_/Q heichips25_sap3/_1316_
+ heichips25_sap3/_1265_ heichips25_sap3__3991_/Q heichips25_sap3/_1317_ heichips25_sap3/net293
+ sg13g2_a221oi_1
XFILLER_3_790 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2961_ net780 VGND VPWR heichips25_can_lehmann_fsm/net1018
+ heichips25_can_lehmann_fsm__2961_/Q clknet_leaf_16_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2892_ net711 VGND VPWR heichips25_can_lehmann_fsm/_0117_
+ heichips25_can_lehmann_fsm__2892_/Q clknet_leaf_18_clk sg13g2_dfrbpq_1
XFILLER_18_0 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1912_ heichips25_can_lehmann_fsm/_1225_ heichips25_can_lehmann_fsm__2931_/Q
+ heichips25_can_lehmann_fsm/net315 VPWR VGND sg13g2_nand2_1
X_08_ uo_out_fsm\[2\] uo_out_sap3\[2\] net507 net37 VPWR VGND sg13g2_mux2_1
Xheichips25_can_lehmann_fsm__1843_ heichips25_can_lehmann_fsm/_1141_ heichips25_can_lehmann_fsm/_1108_
+ heichips25_can_lehmann_fsm/_1157_ heichips25_can_lehmann_fsm/_1159_ VPWR VGND sg13g2_a21o_1
Xheichips25_can_lehmann_fsm__1774_ heichips25_can_lehmann_fsm/_1084_ heichips25_can_lehmann_fsm/_1089_
+ heichips25_can_lehmann_fsm/_1054_ heichips25_can_lehmann_fsm/_1090_ VPWR VGND sg13g2_nand3_1
Xheichips25_can_lehmann_fsm_hold1117 heichips25_can_lehmann_fsm__3056_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1116 sg13g2_dlygate4sd3_1
XFILLER_21_311 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm_hold1128 heichips25_can_lehmann_fsm__3048_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1127 sg13g2_dlygate4sd3_1
XFILLER_33_160 VPWR VGND sg13g2_fill_2
XFILLER_21_333 VPWR VGND sg13g2_fill_2
XFILLER_21_344 VPWR VGND sg13g2_decap_4
XFILLER_22_878 VPWR VGND sg13g2_fill_1
Xheichips25_sap3_hold837 heichips25_sap3/_1256_ VPWR VGND heichips25_sap3/net836 sg13g2_dlygate4sd3_1
XFILLER_21_388 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2326_ heichips25_can_lehmann_fsm/net471 VPWR heichips25_can_lehmann_fsm/_0629_
+ VGND heichips25_can_lehmann_fsm/net933 heichips25_can_lehmann_fsm/net403 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2257_ VGND VPWR heichips25_can_lehmann_fsm/net1183 heichips25_can_lehmann_fsm/net173
+ heichips25_can_lehmann_fsm/_0576_ heichips25_can_lehmann_fsm/_0575_ sg13g2_a21oi_1
Xheichips25_sap3_fanout58 heichips25_sap3/_1052_ heichips25_sap3/net58 VPWR VGND sg13g2_buf_1
Xheichips25_sap3_fanout69 heichips25_sap3/net70 heichips25_sap3/net69 VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm__2188_ VPWR VGND heichips25_can_lehmann_fsm/net164 heichips25_can_lehmann_fsm/_0521_
+ heichips25_can_lehmann_fsm/_0520_ net16 heichips25_can_lehmann_fsm/_0522_ heichips25_can_lehmann_fsm/_0499_
+ sg13g2_a221oi_1
Xoutput38 net38 uo_out[3] VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm__2919__658 VPWR VGND net657 sg13g2_tiehi
Xoutput27 net27 uio_out[0] VPWR VGND sg13g2_buf_1
XFILLER_29_422 VPWR VGND sg13g2_decap_8
XFILLER_17_617 VPWR VGND sg13g2_fill_1
XFILLER_45_959 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2140_ heichips25_sap3/_1496_ heichips25_sap3/_1559_ heichips25_sap3/_1561_
+ VPWR VGND sg13g2_nor2_1
XFILLER_16_138 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__3061__526 VPWR VGND net525 sg13g2_tiehi
XFILLER_40_620 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2071_ heichips25_sap3/_1487_ heichips25_sap3/_1489_ heichips25_sap3/net268
+ heichips25_sap3/_1492_ VPWR VGND sg13g2_nand3_1
XFILLER_25_683 VPWR VGND sg13g2_decap_8
XFILLER_31_119 VPWR VGND sg13g2_fill_2
Xheichips25_sap3_hold1150 heichips25_sap3__4051_/Q VPWR VGND heichips25_sap3/net1149
+ sg13g2_dlygate4sd3_1
XFILLER_12_388 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2973_ heichips25_sap3/_0048_ heichips25_sap3/_0608_ heichips25_sap3/_0609_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__3525_ uio_out_sap3\[5\] heichips25_sap3/net131 heichips25_sap3/_1117_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__3456_ heichips25_sap3/_1060_ heichips25_sap3__3940_/Q heichips25_sap3/net57
+ VPWR VGND sg13g2_nand2_1
XFILLER_48_797 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2407_ heichips25_sap3/_1824_ heichips25_sap3/net80 heichips25_sap3__4024_/Q
+ heichips25_sap3/net86 heichips25_sap3__3952_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__3009__811 VPWR VGND net810 sg13g2_tiehi
XFILLER_47_285 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3387_ heichips25_sap3/_0995_ heichips25_sap3/_0802_ heichips25_sap3/_0872_
+ VPWR VGND sg13g2_xnor2_1
XFILLER_35_458 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2338_ heichips25_sap3/_1486_ heichips25_sap3/_1495_ heichips25_sap3/_1759_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__2269_ heichips25_sap3/_1690_ heichips25_sap3/_1689_ heichips25_sap3/net243
+ heichips25_sap3/_1687_ heichips25_sap3/_1499_ VPWR VGND sg13g2_a22oi_1
XFILLER_15_171 VPWR VGND sg13g2_decap_8
XFILLER_22_119 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__4008_ heichips25_sap3/net445 VGND VPWR heichips25_sap3/_0149_ heichips25_sap3__4008_/Q
+ clkload21/A sg13g2_dfrbpq_1
Xclkbuf_5_25__f_heichips25_sap3\_sap_3_inst.alu_inst.clk heichips25_sap3__4003_/CLK
+ clknet_4_12_0_heichips25_sap3\/sap_3_inst.alu_inst.clk VPWR VGND sg13g2_buf_16
Xclkbuf_0_clk clknet_0_clk clk VPWR VGND sg13g2_buf_16
XFILLER_30_152 VPWR VGND sg13g2_decap_4
XFILLER_7_51 VPWR VGND sg13g2_decap_8
XFILLER_8_871 VPWR VGND sg13g2_fill_2
XFILLER_7_370 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2111_ heichips25_can_lehmann_fsm/_0450_ heichips25_can_lehmann_fsm/net295
+ heichips25_can_lehmann_fsm__2981_/Q heichips25_can_lehmann_fsm/net315 heichips25_can_lehmann_fsm__2933_/Q
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2042_ heichips25_can_lehmann_fsm/net185 VPWR heichips25_can_lehmann_fsm/_0391_
+ VGND heichips25_can_lehmann_fsm/_1074_ heichips25_can_lehmann_fsm/_0390_ sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2944_ net559 VGND VPWR heichips25_can_lehmann_fsm/_0169_
+ heichips25_can_lehmann_fsm__2944_/Q clknet_leaf_22_clk sg13g2_dfrbpq_1
XFILLER_38_241 VPWR VGND sg13g2_decap_8
XFILLER_38_285 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2875_ net745 VGND VPWR heichips25_can_lehmann_fsm/net1016
+ heichips25_can_lehmann_fsm__2875_/Q clknet_leaf_1_clk sg13g2_dfrbpq_1
XFILLER_41_406 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1826_ VPWR heichips25_can_lehmann_fsm/_1142_ heichips25_can_lehmann_fsm/_1141_
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__1757_ heichips25_can_lehmann_fsm/_1077_ heichips25_can_lehmann_fsm/_1074_
+ heichips25_can_lehmann_fsm/_1031_ heichips25_can_lehmann_fsm/_1037_ heichips25_can_lehmann_fsm__2789_/Q
+ VPWR VGND sg13g2_a22oi_1
XFILLER_42_59 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1688_ heichips25_can_lehmann_fsm/_1012_ heichips25_can_lehmann_fsm/net296
+ heichips25_can_lehmann_fsm__2898_/Q heichips25_can_lehmann_fsm/net317 heichips25_can_lehmann_fsm__2994_/Q
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2309_ VGND VPWR heichips25_can_lehmann_fsm/net1188 heichips25_can_lehmann_fsm/net174
+ heichips25_can_lehmann_fsm/_0618_ heichips25_can_lehmann_fsm/_0617_ sg13g2_a21oi_1
Xheichips25_sap3__3310_ heichips25_sap3/_0915_ heichips25_sap3/_0916_ heichips25_sap3/_0919_
+ heichips25_sap3/_0920_ heichips25_sap3/_0921_ VPWR VGND sg13g2_and4_1
XFILLER_18_915 VPWR VGND sg13g2_decap_4
XFILLER_18_959 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3241_ heichips25_sap3/_0841_ heichips25_sap3/_0852_ heichips25_sap3/net61
+ heichips25_sap3/_0854_ VPWR VGND sg13g2_nand3_1
Xheichips25_sap3__3172_ heichips25_sap3/_0785_ heichips25_sap3/_0783_ heichips25_sap3/_0784_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__2123_ heichips25_sap3/_1544_ heichips25_sap3/net236 heichips25_sap3/_1543_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__2054_ VGND VPWR heichips25_sap3/_1475_ heichips25_sap3/_1448_ heichips25_sap3/_1435_
+ sg13g2_or2_1
XFILLER_5_863 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2956_ heichips25_sap3/_0594_ heichips25_sap3/_0590_ heichips25_sap3/_0593_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_can_lehmann_fsm__2937__588 VPWR VGND net587 sg13g2_tiehi
XFILLER_4_362 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2887_ heichips25_sap3/_0520_ heichips25_sap3/_0521_ heichips25_sap3/_0519_
+ heichips25_sap3/_0528_ VPWR VGND heichips25_sap3/_0527_ sg13g2_nand4_1
Xheichips25_sap3__3508_ heichips25_sap3/_1103_ heichips25_sap3/_1101_ heichips25_sap3/_1102_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__3439_ heichips25_sap3/_1045_ heichips25_sap3/net54 heichips25_sap3/_0857_
+ VPWR VGND sg13g2_xnor2_1
XFILLER_35_200 VPWR VGND sg13g2_fill_2
XFILLER_35_244 VPWR VGND sg13g2_fill_1
XFILLER_24_929 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2660_ heichips25_can_lehmann_fsm/net498 VPWR heichips25_can_lehmann_fsm/_0796_
+ VGND heichips25_can_lehmann_fsm/net920 heichips25_can_lehmann_fsm/net384 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__1611_ VPWR heichips25_can_lehmann_fsm/_0935_ heichips25_can_lehmann_fsm/net1056
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__2591_ VGND VPWR heichips25_can_lehmann_fsm/_0900_ heichips25_can_lehmann_fsm/net399
+ heichips25_can_lehmann_fsm/_0195_ heichips25_can_lehmann_fsm/_0761_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__1542_ VPWR heichips25_can_lehmann_fsm/_0866_ heichips25_can_lehmann_fsm/net993
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__2025_ heichips25_can_lehmann_fsm__2781_/Q heichips25_can_lehmann_fsm/net181
+ heichips25_can_lehmann_fsm/_0377_ VPWR VGND sg13g2_nor2_1
X_22__508 VPWR VGND net sg13g2_tielo
XFILLER_37_48 VPWR VGND sg13g2_fill_1
XFILLER_37_37 VPWR VGND sg13g2_decap_8
XFILLER_27_745 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2927_ net627 VGND VPWR heichips25_can_lehmann_fsm/_0152_
+ heichips25_can_lehmann_fsm__2927_/Q clknet_leaf_13_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2858_ net779 VGND VPWR heichips25_can_lehmann_fsm/_0083_
+ heichips25_can_lehmann_fsm__2858_/Q clknet_leaf_10_clk sg13g2_dfrbpq_1
XFILLER_26_255 VPWR VGND sg13g2_fill_1
XFILLER_27_767 VPWR VGND sg13g2_fill_1
XFILLER_14_417 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1809_ VGND VPWR heichips25_can_lehmann_fsm__2899_/Q heichips25_can_lehmann_fsm/net296
+ heichips25_can_lehmann_fsm/_1125_ heichips25_can_lehmann_fsm/net300 sg13g2_a21oi_1
XFILLER_26_299 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2789_ net628 VGND VPWR heichips25_can_lehmann_fsm/net1247
+ heichips25_can_lehmann_fsm__2789_/Q clknet_leaf_1_clk sg13g2_dfrbpq_1
Xheichips25_sap3__2810_ VGND VPWR heichips25_sap3/_0455_ heichips25_sap3/_0454_ heichips25_sap3/net204
+ sg13g2_or2_1
Xheichips25_sap3__3790_ heichips25_sap3/_1296_ heichips25_sap3/_1298_ heichips25_sap3/_1295_
+ heichips25_sap3/_1300_ VPWR VGND heichips25_sap3/_1299_ sg13g2_nand4_1
Xheichips25_can_lehmann_fsm__2973__733 VPWR VGND net732 sg13g2_tiehi
Xheichips25_sap3__2741_ heichips25_sap3/_0387_ heichips25_sap3/net283 heichips25_sap3__3918_/Q
+ VPWR VGND sg13g2_nand2b_1
Xheichips25_sap3__2672_ heichips25_sap3/_1593_ heichips25_sap3/_1803_ heichips25_sap3/_1811_
+ uio_oe_sap3\[6\] VPWR VGND sg13g2_nor3_1
XFILLER_49_303 VPWR VGND sg13g2_fill_1
XFILLER_49_347 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3224_ heichips25_sap3/net152 heichips25_sap3/_0762_ heichips25_sap3__3949_/Q
+ heichips25_sap3/_0837_ VPWR VGND sg13g2_nand3_1
Xheichips25_sap3__3155_ heichips25_sap3/_0666_ heichips25_sap3/_0678_ heichips25_sap3/_0697_
+ heichips25_sap3/_0768_ VPWR VGND sg13g2_nor3_1
XFILLER_32_247 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3086_ heichips25_sap3/_1525_ heichips25_sap3/_1535_ heichips25_sap3/_0638_
+ heichips25_sap3/_0698_ heichips25_sap3/_0699_ VPWR VGND sg13g2_nor4_1
Xheichips25_sap3__2106_ heichips25_sap3/_1436_ heichips25_sap3/_1489_ heichips25_sap3/_1434_
+ heichips25_sap3/_1527_ VPWR VGND sg13g2_nand3_1
XFILLER_32_269 VPWR VGND sg13g2_decap_8
XFILLER_13_494 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2037_ VGND VPWR heichips25_sap3/_1458_ heichips25_sap3/net250 heichips25_sap3/net251
+ sg13g2_or2_1
XFILLER_9_454 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3988_ heichips25_sap3/net443 VGND VPWR heichips25_sap3/_0129_ heichips25_sap3__3988_/Q
+ heichips25_sap3__3988_/CLK sg13g2_dfrbpq_1
Xheichips25_sap3__2939_ heichips25_sap3/_0553_ heichips25_sap3/_0577_ heichips25_sap3/_0578_
+ VPWR VGND sg13g2_and2_1
XFILLER_28_509 VPWR VGND sg13g2_fill_1
XFILLER_48_380 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2712_ heichips25_can_lehmann_fsm/net485 VPWR heichips25_can_lehmann_fsm/_0822_
+ VGND heichips25_can_lehmann_fsm__3031_/Q heichips25_can_lehmann_fsm/net417 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2643_ VGND VPWR heichips25_can_lehmann_fsm/_0887_ heichips25_can_lehmann_fsm/net399
+ heichips25_can_lehmann_fsm/_0221_ heichips25_can_lehmann_fsm/_0787_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2574_ heichips25_can_lehmann_fsm/net482 VPWR heichips25_can_lehmann_fsm/_0753_
+ VGND heichips25_can_lehmann_fsm/net1038 heichips25_can_lehmann_fsm/net409 sg13g2_o21ai_1
XFILLER_20_910 VPWR VGND sg13g2_fill_2
XFILLER_23_28 VPWR VGND sg13g2_decap_8
XFILLER_20_943 VPWR VGND sg13g2_fill_1
XFILLER_23_39 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__3057_ net557 VGND VPWR heichips25_can_lehmann_fsm/_0282_
+ heichips25_can_lehmann_fsm__3057_/Q clknet_leaf_16_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2008_ heichips25_can_lehmann_fsm__2787_/Q VPWR heichips25_can_lehmann_fsm/_0362_
+ VGND heichips25_can_lehmann_fsm__2786_/Q heichips25_can_lehmann_fsm/_1068_ sg13g2_o21ai_1
Xclkbuf_4_13_0_heichips25_sap3\_sap_3_inst.alu_inst.clk clknet_0_heichips25_sap3\/sap_3_inst.alu_inst.clk
+ clknet_4_13_0_heichips25_sap3\/sap_3_inst.alu_inst.clk VPWR VGND sg13g2_buf_8
XFILLER_27_586 VPWR VGND sg13g2_fill_2
XFILLER_14_225 VPWR VGND sg13g2_fill_1
XFILLER_14_236 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3911_ heichips25_sap3/net455 VGND VPWR heichips25_sap3/_0052_ heichips25_sap3__3911_/Q
+ clkload25/A sg13g2_dfrbpq_1
XFILLER_11_987 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3842_ heichips25_sap3/net1224 VPWR heichips25_sap3/_1344_ VGND heichips25_sap3/_0018_
+ heichips25_sap3/_1260_ sg13g2_o21ai_1
XFILLER_7_969 VPWR VGND sg13g2_fill_1
XFILLER_6_479 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3773_ VGND VPWR heichips25_sap3/_1392_ heichips25_sap3/net290 heichips25_sap3/_1285_
+ heichips25_sap3/net339 sg13g2_a21oi_1
Xheichips25_sap3__2724_ VGND VPWR heichips25_sap3/_0350_ heichips25_sap3/_0369_ heichips25_sap3/_0370_
+ heichips25_sap3/_0349_ sg13g2_a21oi_1
XFILLER_2_663 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2655_ VGND VPWR heichips25_sap3/_0318_ heichips25_sap3/_0320_ heichips25_sap3/_0322_
+ heichips25_sap3/_1455_ sg13g2_a21oi_1
Xheichips25_sap3__2586_ heichips25_sap3/net284 heichips25_sap3/net156 heichips25_sap3/_0259_
+ VPWR VGND sg13g2_nor2_1
XFILLER_18_531 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3207_ heichips25_sap3/_0816_ heichips25_sap3/_0817_ heichips25_sap3/_0815_
+ heichips25_sap3/_0820_ VPWR VGND heichips25_sap3/_0818_ sg13g2_nand4_1
Xheichips25_sap3__3138_ heichips25_sap3/_0667_ heichips25_sap3/_0679_ heichips25_sap3/_0751_
+ VPWR VGND sg13g2_nor2_1
XFILLER_33_589 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2802__603 VPWR VGND net602 sg13g2_tiehi
Xheichips25_sap3__3069_ heichips25_sap3/_0682_ heichips25_sap3/_0681_ heichips25_sap3/_1486_
+ heichips25_sap3/_1754_ heichips25_sap3/_1685_ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2290_ VGND VPWR heichips25_can_lehmann_fsm/net207 heichips25_can_lehmann_fsm/_0601_
+ heichips25_can_lehmann_fsm/_0053_ heichips25_can_lehmann_fsm/_0602_ sg13g2_a21oi_1
Xclkload10 VPWR clkload10/Y clknet_leaf_16_clk VGND sg13g2_inv_1
Xclkload21 VPWR clkload21/Y clkload21/A VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm_fanout305 heichips25_can_lehmann_fsm/net309 heichips25_can_lehmann_fsm/net305
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout327 heichips25_can_lehmann_fsm/net329 heichips25_can_lehmann_fsm/net327
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout338 heichips25_can_lehmann_fsm/_0983_ heichips25_can_lehmann_fsm/net338
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout316 heichips25_can_lehmann_fsm/_0993_ heichips25_can_lehmann_fsm/net316
+ VPWR VGND sg13g2_buf_1
XFILLER_47_1027 VPWR VGND sg13g2_fill_2
XFILLER_47_1016 VPWR VGND sg13g2_decap_8
XFILLER_48_0 VPWR VGND sg13g2_decap_4
XFILLER_5_490 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_fanout349 heichips25_can_lehmann_fsm/net350 heichips25_can_lehmann_fsm/net349
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm__2852__792 VPWR VGND net791 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2626_ heichips25_can_lehmann_fsm/net478 VPWR heichips25_can_lehmann_fsm/_0779_
+ VGND heichips25_can_lehmann_fsm/net963 heichips25_can_lehmann_fsm/net409 sg13g2_o21ai_1
XFILLER_24_567 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2557_ VGND VPWR heichips25_can_lehmann_fsm/_0908_ heichips25_can_lehmann_fsm/net382
+ heichips25_can_lehmann_fsm/_0178_ heichips25_can_lehmann_fsm/_0744_ sg13g2_a21oi_1
Xclkload4 clkload4/Y clknet_leaf_2_clk VPWR VGND sg13g2_inv_2
Xheichips25_can_lehmann_fsm__2488_ heichips25_can_lehmann_fsm/net464 VPWR heichips25_can_lehmann_fsm/_0710_
+ VGND heichips25_can_lehmann_fsm/net1070 heichips25_can_lehmann_fsm/net358 sg13g2_o21ai_1
X_28__514 VPWR VGND net513 sg13g2_tielo
Xheichips25_sap3__2440_ heichips25_sap3/_1855_ heichips25_sap3/net156 heichips25_sap3/_1854_
+ VPWR VGND sg13g2_nand2_1
XFILLER_47_637 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2371_ heichips25_sap3/_1792_ heichips25_sap3/_1771_ heichips25_sap3/_1791_
+ VPWR VGND sg13g2_nand2_1
XFILLER_15_501 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__4041_ heichips25_sap3/net460 VGND VPWR heichips25_sap3/net1179 heichips25_sap3__4041_/Q
+ clknet_leaf_3_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2784__639 VPWR VGND net638 sg13g2_tiehi
XFILLER_15_534 VPWR VGND sg13g2_fill_1
XFILLER_43_865 VPWR VGND sg13g2_fill_1
XFILLER_42_375 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm_hold950 heichips25_can_lehmann_fsm/_0086_ VPWR VGND heichips25_can_lehmann_fsm/net949
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold961 heichips25_can_lehmann_fsm__3026_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net960 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold983 heichips25_can_lehmann_fsm/_0145_ VPWR VGND heichips25_can_lehmann_fsm/net982
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold972 heichips25_can_lehmann_fsm/_0167_ VPWR VGND heichips25_can_lehmann_fsm/net971
+ sg13g2_dlygate4sd3_1
XFILLER_11_773 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm_hold994 heichips25_can_lehmann_fsm__3032_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net993 sg13g2_dlygate4sd3_1
XFILLER_10_294 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3825_ heichips25_sap3/_1331_ heichips25_sap3/_1265_ heichips25_sap3__4001_/Q
+ heichips25_sap3/net293 heichips25_sap3__3993_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_6_298 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3756_ heichips25_sap3/_1268_ heichips25_sap3/net292 heichips25_sap3__3955_/Q
+ heichips25_sap3/_1265_ heichips25_sap3__3995_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2707_ heichips25_sap3/net278 heichips25_sap3__3920_/Q heichips25_sap3/_0353_
+ VPWR VGND sg13g2_nor2_1
XFILLER_34_6 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3687_ heichips25_sap3/_1225_ heichips25_sap3__4006_/Q heichips25_sap3/net113
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__2638_ VGND VPWR heichips25_sap3/net235 heichips25_sap3/_1560_ heichips25_sap3/_0305_
+ heichips25_sap3/_1558_ sg13g2_a21oi_1
XFILLER_37_114 VPWR VGND sg13g2_decap_8
XFILLER_37_103 VPWR VGND sg13g2_fill_2
XFILLER_37_147 VPWR VGND sg13g2_decap_4
XFILLER_37_125 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2569_ VGND VPWR heichips25_sap3/_0243_ heichips25_sap3/_0214_ heichips25_sap3/_1878_
+ sg13g2_or2_1
X_24_ net509 uio_oe_sap3\[2\] net505 net21 VPWR VGND sg13g2_mux2_1
Xheichips25_can_lehmann_fsm__1790_ heichips25_can_lehmann_fsm__2816_/Q heichips25_can_lehmann_fsm/_1105_
+ heichips25_can_lehmann_fsm/_1106_ VPWR VGND sg13g2_nor2b_1
XFILLER_37_169 VPWR VGND sg13g2_decap_4
XFILLER_1_97 VPWR VGND sg13g2_fill_1
XFILLER_19_884 VPWR VGND sg13g2_fill_1
XFILLER_46_692 VPWR VGND sg13g2_fill_2
XFILLER_34_843 VPWR VGND sg13g2_fill_2
XFILLER_34_832 VPWR VGND sg13g2_decap_8
XFILLER_18_394 VPWR VGND sg13g2_decap_8
XFILLER_19_895 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2411_ VGND VPWR heichips25_can_lehmann_fsm/_0947_ heichips25_can_lehmann_fsm/net421
+ heichips25_can_lehmann_fsm/_0105_ heichips25_can_lehmann_fsm/_0671_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2342_ heichips25_can_lehmann_fsm/net494 VPWR heichips25_can_lehmann_fsm/_0637_
+ VGND heichips25_can_lehmann_fsm/net1034 heichips25_can_lehmann_fsm/net406 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2273_ VGND VPWR heichips25_can_lehmann_fsm/net965 heichips25_can_lehmann_fsm/net172
+ heichips25_can_lehmann_fsm/_0589_ heichips25_can_lehmann_fsm/_0588_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm_fanout179 heichips25_can_lehmann_fsm/net180 heichips25_can_lehmann_fsm/net179
+ VPWR VGND sg13g2_buf_1
XFILLER_29_27 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1988_ VGND VPWR heichips25_can_lehmann_fsm/net177 heichips25_can_lehmann_fsm/_0344_
+ heichips25_can_lehmann_fsm/_0008_ heichips25_can_lehmann_fsm/_0345_ sg13g2_a21oi_1
XFILLER_12_548 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2609_ VGND VPWR heichips25_can_lehmann_fsm/_0895_ heichips25_can_lehmann_fsm/net381
+ heichips25_can_lehmann_fsm/_0204_ heichips25_can_lehmann_fsm/_0770_ sg13g2_a21oi_1
Xheichips25_sap3__1940_ VPWR heichips25_sap3/_1366_ heichips25_sap3/net830 VGND sg13g2_inv_1
XFILLER_3_202 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3610_ heichips25_sap3/_1141_ heichips25_sap3__3977_/Q heichips25_sap3/_1171_
+ heichips25_sap3/_0118_ VPWR VGND sg13g2_mux2_1
Xheichips25_sap3__3541_ VGND VPWR heichips25_sap3/_1042_ heichips25_sap3/_1043_ heichips25_sap3/_1131_
+ heichips25_sap3/net120 sg13g2_a21oi_1
XFILLER_0_964 VPWR VGND sg13g2_decap_8
XFILLER_48_946 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3472_ heichips25_sap3/net57 heichips25_sap3__3943_/Q heichips25_sap3/_1072_
+ heichips25_sap3/_0084_ VPWR VGND sg13g2_a21o_1
XFILLER_19_103 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2423_ VPWR VGND heichips25_sap3__4008_/Q heichips25_sap3/net80 heichips25_sap3/net74
+ heichips25_sap3__4016_/Q heichips25_sap3/_1840_ heichips25_sap3/net217 sg13g2_a221oi_1
Xheichips25_sap3__2354_ VGND VPWR heichips25_sap3/_1775_ heichips25_sap3/_1774_ heichips25_sap3/net266
+ sg13g2_or2_1
XFILLER_19_158 VPWR VGND sg13g2_decap_4
XFILLER_16_821 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__4024_ heichips25_sap3/net442 VGND VPWR heichips25_sap3/_0165_ heichips25_sap3__4024_/Q
+ heichips25_sap3__4024_/CLK sg13g2_dfrbpq_1
Xheichips25_sap3__2285_ heichips25_sap3/net223 VPWR heichips25_sap3/_1706_ VGND heichips25_sap3/_1701_
+ heichips25_sap3/_1703_ sg13g2_o21ai_1
XFILLER_16_865 VPWR VGND sg13g2_decap_4
XFILLER_37_1026 VPWR VGND sg13g2_fill_2
XFILLER_15_364 VPWR VGND sg13g2_decap_4
XFILLER_15_386 VPWR VGND sg13g2_fill_1
XFILLER_30_301 VPWR VGND sg13g2_fill_2
XFILLER_30_389 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3808_ heichips25_sap3/_1313_ heichips25_sap3/_1314_ heichips25_sap3/_1312_
+ heichips25_sap3/_1316_ VPWR VGND heichips25_sap3/_1315_ sg13g2_nand4_1
Xheichips25_sap3__3739_ heichips25_sap3/net1130 heichips25_sap3/net1176 heichips25_sap3/_1254_
+ VPWR VGND sg13g2_nor2_1
XFILLER_39_913 VPWR VGND sg13g2_fill_1
XFILLER_38_401 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2960_ net784 VGND VPWR heichips25_can_lehmann_fsm/net1046
+ heichips25_can_lehmann_fsm__2960_/Q clknet_leaf_16_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2891_ net713 VGND VPWR heichips25_can_lehmann_fsm/net956
+ heichips25_can_lehmann_fsm__2891_/Q clknet_leaf_18_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1911_ VGND VPWR heichips25_can_lehmann_fsm__3051_/Q heichips25_can_lehmann_fsm/_1161_
+ heichips25_can_lehmann_fsm/_1224_ heichips25_can_lehmann_fsm/_1139_ sg13g2_a21oi_1
X_07_ uo_out_fsm\[1\] uo_out_sap3\[1\] net504 net36 VPWR VGND sg13g2_mux2_1
Xheichips25_can_lehmann_fsm__1842_ heichips25_can_lehmann_fsm/_1153_ heichips25_can_lehmann_fsm__3060_/Q
+ heichips25_can_lehmann_fsm/_1157_ heichips25_can_lehmann_fsm/_1158_ VPWR VGND sg13g2_a21o_1
XFILLER_26_629 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1773_ heichips25_can_lehmann_fsm/_1086_ heichips25_can_lehmann_fsm/_1087_
+ heichips25_can_lehmann_fsm/_1085_ heichips25_can_lehmann_fsm/_1089_ VPWR VGND heichips25_can_lehmann_fsm/_1088_
+ sg13g2_nand4_1
XFILLER_25_139 VPWR VGND sg13g2_fill_2
XFILLER_15_18 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm_hold1107 heichips25_can_lehmann_fsm__2935_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1106 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1118 heichips25_can_lehmann_fsm__3049_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1117 sg13g2_dlygate4sd3_1
XFILLER_22_846 VPWR VGND sg13g2_decap_4
XFILLER_22_868 VPWR VGND sg13g2_decap_4
Xheichips25_sap3_hold838 heichips25_sap3/_0172_ VPWR VGND heichips25_sap3/net837 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__2325_ VGND VPWR heichips25_can_lehmann_fsm/_0970_ heichips25_can_lehmann_fsm/net363
+ heichips25_can_lehmann_fsm/_0062_ heichips25_can_lehmann_fsm/_0628_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2256_ heichips25_can_lehmann_fsm/net173 heichips25_can_lehmann_fsm/_0574_
+ heichips25_can_lehmann_fsm/_0575_ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3_fanout59 heichips25_sap3/_0830_ heichips25_sap3/net59 VPWR VGND sg13g2_buf_1
Xheichips25_sap3_fanout48 heichips25_sap3/net49 heichips25_sap3/net48 VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm__2187_ heichips25_can_lehmann_fsm/_0969_ heichips25_can_lehmann_fsm/_0494_
+ heichips25_can_lehmann_fsm/_0521_ VPWR VGND sg13g2_nor2_1
Xoutput39 net39 uo_out[4] VPWR VGND sg13g2_buf_1
Xoutput28 net28 uio_out[1] VPWR VGND sg13g2_buf_1
XFILLER_0_227 VPWR VGND sg13g2_fill_2
XFILLER_5_1024 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2070_ heichips25_sap3/net257 heichips25_sap3/net255 heichips25_sap3/_1490_
+ heichips25_sap3/_1491_ VPWR VGND sg13g2_nor3_1
XFILLER_12_356 VPWR VGND sg13g2_fill_2
Xclkbuf_5_8__f_heichips25_sap3\_sap_3_inst.alu_inst.clk heichips25_sap3__4017_/CLK
+ clknet_4_4_0_heichips25_sap3\/sap_3_inst.alu_inst.clk VPWR VGND sg13g2_buf_16
Xheichips25_sap3__2972_ heichips25_sap3/_0609_ heichips25_sap3/net153 heichips25_sap3/_0372_
+ heichips25_sap3/net167 heichips25_sap3__3899_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_4_544 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3524_ heichips25_sap3/net120 heichips25_sap3/_1001_ heichips25_sap3/_1116_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__3455_ VPWR heichips25_sap3/_0080_ heichips25_sap3/_1059_ VGND sg13g2_inv_1
Xheichips25_sap3__2406_ heichips25_sap3__3896_/Q net43 heichips25_sap3/net215 heichips25_sap3/_0037_
+ VPWR VGND sg13g2_mux2_1
Xheichips25_sap3__3386_ heichips25_sap3/_0994_ heichips25_sap3/_0970_ heichips25_sap3/_0991_
+ VPWR VGND sg13g2_xnor2_1
Xheichips25_sap3__2337_ heichips25_sap3/_1758_ heichips25_sap3/net245 heichips25_sap3/_1757_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__2268_ heichips25_sap3/net229 heichips25_sap3/_1553_ heichips25_sap3/net235
+ heichips25_sap3/_1689_ VPWR VGND heichips25_sap3/_1681_ sg13g2_nand4_1
XFILLER_31_610 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__4007_ heichips25_sap3/net445 VGND VPWR heichips25_sap3/_0148_ heichips25_sap3__4007_/Q
+ clkload21/A sg13g2_dfrbpq_1
Xheichips25_sap3__2199_ heichips25_sap3/_1448_ heichips25_sap3/_1615_ heichips25_sap3/_1620_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_can_lehmann_fsm__2110_ heichips25_can_lehmann_fsm/_0449_ heichips25_can_lehmann_fsm/net298
+ heichips25_can_lehmann_fsm__2909_/Q heichips25_can_lehmann_fsm/net308 heichips25_can_lehmann_fsm__2957_/Q
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2041_ VGND VPWR heichips25_can_lehmann_fsm/_0979_ heichips25_can_lehmann_fsm/_1073_
+ heichips25_can_lehmann_fsm/_0390_ heichips25_can_lehmann_fsm/_0978_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2943_ net563 VGND VPWR heichips25_can_lehmann_fsm/net1026
+ heichips25_can_lehmann_fsm__2943_/Q clknet_leaf_22_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2874_ net747 VGND VPWR heichips25_can_lehmann_fsm/_0099_
+ heichips25_can_lehmann_fsm__2874_/Q clknet_leaf_0_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2810__587 VPWR VGND net586 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__1825_ heichips25_can_lehmann_fsm__3045_/Q heichips25_can_lehmann_fsm__3044_/Q
+ heichips25_can_lehmann_fsm/net343 heichips25_can_lehmann_fsm/_1141_ VPWR VGND sg13g2_nor3_1
Xheichips25_can_lehmann_fsm__1756_ heichips25_can_lehmann_fsm/_1076_ heichips25_can_lehmann_fsm/net345
+ heichips25_can_lehmann_fsm/_1032_ VPWR VGND sg13g2_nand2_1
Xheichips25_can_lehmann_fsm__1687_ VGND VPWR heichips25_can_lehmann_fsm__2946_/Q heichips25_can_lehmann_fsm/net305
+ heichips25_can_lehmann_fsm/_1011_ heichips25_can_lehmann_fsm/net300 sg13g2_a21oi_1
XFILLER_22_654 VPWR VGND sg13g2_fill_1
XFILLER_21_197 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2308_ heichips25_can_lehmann_fsm/net174 heichips25_can_lehmann_fsm/_0616_
+ heichips25_can_lehmann_fsm/_0617_ VPWR VGND sg13g2_nor2_1
Xheichips25_can_lehmann_fsm__2239_ heichips25_can_lehmann_fsm__2818_/Q heichips25_can_lehmann_fsm/net1174
+ heichips25_can_lehmann_fsm/_0561_ VPWR VGND sg13g2_xor2_1
XFILLER_49_518 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3240_ heichips25_sap3/_0853_ heichips25_sap3/_0841_ heichips25_sap3/_0852_
+ VPWR VGND sg13g2_nand2_1
XFILLER_17_415 VPWR VGND sg13g2_fill_2
XFILLER_45_757 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3171_ heichips25_sap3/_0784_ heichips25_sap3/net144 heichips25_sap3__3970_/Q
+ heichips25_sap3/net128 heichips25_sap3__3946_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2122_ heichips25_sap3/_1543_ heichips25_sap3/net265 heichips25_sap3/_1542_
+ VPWR VGND sg13g2_xnor2_1
XFILLER_25_470 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2053_ heichips25_sap3/_1435_ heichips25_sap3/_1448_ heichips25_sap3/_1474_
+ VPWR VGND sg13g2_nor2_1
XFILLER_13_621 VPWR VGND sg13g2_fill_1
XFILLER_13_643 VPWR VGND sg13g2_fill_2
XFILLER_40_462 VPWR VGND sg13g2_fill_1
XFILLER_12_131 VPWR VGND sg13g2_fill_2
XFILLER_40_484 VPWR VGND sg13g2_decap_4
XFILLER_8_179 VPWR VGND sg13g2_fill_1
XFILLER_8_168 VPWR VGND sg13g2_decap_8
XFILLER_5_842 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2955_ heichips25_sap3/_0593_ heichips25_sap3/_1895_ heichips25_sap3/_0347_
+ VPWR VGND sg13g2_nand2b_1
XFILLER_4_352 VPWR VGND sg13g2_fill_1
XFILLER_4_385 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2886_ VPWR VGND heichips25_sap3/_0340_ heichips25_sap3/_0526_ heichips25_sap3/_0524_
+ heichips25_sap3/_0338_ heichips25_sap3/_0527_ heichips25_sap3/_0523_ sg13g2_a221oi_1
Xheichips25_sap3__3507_ VGND VPWR uio_oe_sap3\[2\] heichips25_sap3/_1087_ heichips25_sap3/_1102_
+ heichips25_sap3/net122 sg13g2_a21oi_1
Xheichips25_sap3__3438_ heichips25_sap3/_1042_ heichips25_sap3/_1043_ heichips25_sap3/net125
+ heichips25_sap3/_1044_ VPWR VGND sg13g2_nand3_1
Xheichips25_sap3__3369_ heichips25_sap3/_0978_ heichips25_sap3/net63 heichips25_sap3/_0855_
+ VPWR VGND sg13g2_xnor2_1
XFILLER_35_278 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2590_ heichips25_can_lehmann_fsm/net480 VPWR heichips25_can_lehmann_fsm/_0761_
+ VGND heichips25_can_lehmann_fsm__2970_/Q heichips25_can_lehmann_fsm/net399 sg13g2_o21ai_1
XFILLER_23_429 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__1610_ VPWR heichips25_can_lehmann_fsm/_0934_ heichips25_can_lehmann_fsm/net1008
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__1541_ VPWR heichips25_can_lehmann_fsm/_0865_ heichips25_can_lehmann_fsm/net1160
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__2024_ heichips25_can_lehmann_fsm/_0376_ heichips25_can_lehmann_fsm/net184
+ heichips25_can_lehmann_fsm/_0374_ heichips25_can_lehmann_fsm/net197 heichips25_can_lehmann_fsm__2788_/Q
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2926_ net631 VGND VPWR heichips25_can_lehmann_fsm/net1048
+ heichips25_can_lehmann_fsm__2926_/Q clknet_leaf_13_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2857_ net781 VGND VPWR heichips25_can_lehmann_fsm/_0082_
+ heichips25_can_lehmann_fsm__2857_/Q clknet_leaf_10_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1808_ heichips25_can_lehmann_fsm/_1124_ heichips25_can_lehmann_fsm/net331
+ heichips25_can_lehmann_fsm/net343 heichips25_can_lehmann_fsm/net313 heichips25_can_lehmann_fsm__2923_/Q
+ VPWR VGND sg13g2_a22oi_1
XFILLER_42_749 VPWR VGND sg13g2_fill_1
XFILLER_23_941 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2788_ net630 VGND VPWR heichips25_can_lehmann_fsm/_0013_
+ heichips25_can_lehmann_fsm__2788_/Q clknet_leaf_1_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1739_ VGND VPWR heichips25_can_lehmann_fsm/_1059_ heichips25_can_lehmann_fsm/net344
+ heichips25_can_lehmann_fsm__2801_/Q sg13g2_or2_1
Xheichips25_can_lehmann_fsm__2862__772 VPWR VGND net771 sg13g2_tiehi
XFILLER_10_613 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2740_ heichips25_sap3/_0386_ heichips25_sap3/net279 heichips25_sap3__3920_/Q
+ VPWR VGND sg13g2_nand2b_1
Xheichips25_sap3__2671_ VPWR VGND heichips25_sap3/_1827_ heichips25_sap3/net66 heichips25_sap3/_1830_
+ heichips25_sap3/_1404_ uio_oe_sap3\[5\] heichips25_sap3/net91 sg13g2_a221oi_1
XFILLER_17_212 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3223_ heichips25_sap3/net152 heichips25_sap3/net150 heichips25_sap3__3957_/Q
+ heichips25_sap3/_0836_ VPWR VGND sg13g2_nand3_1
XFILLER_17_256 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3154_ heichips25_sap3/_0767_ heichips25_sap3/_0696_ heichips25_sap3/net150
+ VPWR VGND sg13g2_nand2_1
Xclkbuf_2_0__f_clk clknet_2_0__leaf_clk clknet_0_clk VPWR VGND sg13g2_buf_16
Xheichips25_can_lehmann_fsm__2980__705 VPWR VGND net704 sg13g2_tiehi
XFILLER_33_705 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2105_ heichips25_sap3/_1435_ heichips25_sap3/_1437_ heichips25_sap3/_1490_
+ heichips25_sap3/_1526_ VPWR VGND sg13g2_nor3_1
Xheichips25_sap3__3085_ heichips25_sap3/_0297_ VPWR heichips25_sap3/_0698_ VGND heichips25_sap3/_1495_
+ heichips25_sap3/_1625_ sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2908__680 VPWR VGND net679 sg13g2_tiehi
XFILLER_9_422 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2036_ heichips25_sap3/net251 heichips25_sap3/net250 heichips25_sap3/_1457_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_can_lehmann_fsm__2794__619 VPWR VGND net618 sg13g2_tiehi
Xheichips25_sap3__3987_ heichips25_sap3/net457 VGND VPWR heichips25_sap3/_0128_ heichips25_sap3__3987_/Q
+ heichips25_sap3__3990_/CLK sg13g2_dfrbpq_1
Xheichips25_sap3__2938_ heichips25_sap3/_0552_ VPWR heichips25_sap3/_0577_ VGND heichips25_sap3/net279
+ heichips25_sap3/net211 sg13g2_o21ai_1
XFILLER_4_160 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2869_ heichips25_sap3/_0499_ heichips25_sap3/_0508_ heichips25_sap3/_0509_
+ heichips25_sap3/_0510_ heichips25_sap3/_0511_ VPWR VGND sg13g2_and4_1
XFILLER_4_53 VPWR VGND sg13g2_decap_8
XFILLER_36_554 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2711_ VGND VPWR heichips25_can_lehmann_fsm/_0867_ heichips25_can_lehmann_fsm/net378
+ heichips25_can_lehmann_fsm/_0255_ heichips25_can_lehmann_fsm/_0821_ sg13g2_a21oi_1
Xclkbuf_5_26__f_heichips25_sap3\_sap_3_inst.alu_inst.clk heichips25_sap3__4021_/CLK
+ clknet_4_13_0_heichips25_sap3\/sap_3_inst.alu_inst.clk VPWR VGND sg13g2_buf_16
Xheichips25_can_lehmann_fsm__2642_ heichips25_can_lehmann_fsm/net469 VPWR heichips25_can_lehmann_fsm/_0787_
+ VGND heichips25_can_lehmann_fsm/net1090 heichips25_can_lehmann_fsm/net399 sg13g2_o21ai_1
XFILLER_23_226 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2573_ VGND VPWR heichips25_can_lehmann_fsm/_0904_ heichips25_can_lehmann_fsm/net374
+ heichips25_can_lehmann_fsm/_0186_ heichips25_can_lehmann_fsm/_0752_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__3056_ net621 VGND VPWR heichips25_can_lehmann_fsm/_0281_
+ heichips25_can_lehmann_fsm__3056_/Q clknet_leaf_16_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2007_ VPWR VGND heichips25_can_lehmann_fsm/net191 heichips25_can_lehmann_fsm/_0361_
+ heichips25_can_lehmann_fsm/_0360_ heichips25_can_lehmann_fsm/_0357_ heichips25_can_lehmann_fsm/_0011_
+ heichips25_can_lehmann_fsm/_0359_ sg13g2_a221oi_1
Xheichips25_can_lehmann_fsm__2909_ net677 VGND VPWR heichips25_can_lehmann_fsm/_0134_
+ heichips25_can_lehmann_fsm__2909_/Q clknet_leaf_15_clk sg13g2_dfrbpq_1
XFILLER_27_532 VPWR VGND sg13g2_decap_8
XFILLER_14_204 VPWR VGND sg13g2_decap_8
XFILLER_11_900 VPWR VGND sg13g2_decap_4
XFILLER_14_259 VPWR VGND sg13g2_decap_4
XFILLER_22_270 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3910_ heichips25_sap3/net448 VGND VPWR heichips25_sap3/_0051_ heichips25_sap3__3910_/Q
+ clkload24/A sg13g2_dfrbpq_1
XFILLER_10_487 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3841_ heichips25_sap3/_1343_ heichips25_sap3/net1178 heichips25_sap3/_0182_
+ VPWR VGND sg13g2_xor2_1
XFILLER_13_95 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3772_ heichips25_sap3/_1277_ heichips25_sap3/_1280_ heichips25_sap3/_1273_
+ heichips25_sap3/_1284_ VPWR VGND heichips25_sap3/_1283_ sg13g2_nand4_1
Xheichips25_sap3__2723_ VGND VPWR heichips25_sap3/_0352_ heichips25_sap3/_0368_ heichips25_sap3/_0369_
+ heichips25_sap3/_0353_ sg13g2_a21oi_1
XFILLER_49_123 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2654_ heichips25_sap3/net227 VPWR heichips25_sap3/_0321_ VGND heichips25_sap3/net249
+ heichips25_sap3/net248 sg13g2_o21ai_1
XFILLER_1_174 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2585_ net5 heichips25_sap3/_1770_ heichips25_sap3/_0258_ VPWR VGND
+ sg13g2_and2_1
XFILLER_46_896 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3206_ heichips25_sap3/_0815_ heichips25_sap3/_0816_ heichips25_sap3/_0817_
+ heichips25_sap3/_0818_ heichips25_sap3/_0819_ VPWR VGND sg13g2_and4_1
XFILLER_33_513 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3137_ heichips25_sap3/_0750_ heichips25_sap3/_0731_ heichips25_sap3/net166
+ VPWR VGND sg13g2_nand2_1
XFILLER_33_579 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3068_ heichips25_sap3/_1526_ heichips25_sap3/_1568_ heichips25_sap3/_1507_
+ heichips25_sap3/_0681_ VPWR VGND sg13g2_nand3_1
Xheichips25_sap3__2019_ heichips25_sap3/_1435_ heichips25_sap3/_1437_ heichips25_sap3/_1438_
+ heichips25_sap3/_1439_ heichips25_sap3/_1440_ VPWR VGND sg13g2_nor4_1
Xclkload22 VPWR clkload22/Y clkload22/A VGND sg13g2_inv_1
Xclkload11 clknet_leaf_17_clk clkload11/X VPWR VGND sg13g2_buf_8
Xheichips25_can_lehmann_fsm_fanout328 heichips25_can_lehmann_fsm/net330 heichips25_can_lehmann_fsm/net328
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout306 heichips25_can_lehmann_fsm/net309 heichips25_can_lehmann_fsm/net306
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout317 heichips25_can_lehmann_fsm/net320 heichips25_can_lehmann_fsm/net317
+ VPWR VGND sg13g2_buf_1
Xheichips25_sap3__2003__815 VPWR net814 heichips25_sap3__4005_/CLK VGND sg13g2_inv_1
XFILLER_24_546 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2625_ VGND VPWR heichips25_can_lehmann_fsm/_0891_ heichips25_can_lehmann_fsm/net374
+ heichips25_can_lehmann_fsm/_0212_ heichips25_can_lehmann_fsm/_0778_ sg13g2_a21oi_1
XFILLER_12_708 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2556_ heichips25_can_lehmann_fsm/net495 VPWR heichips25_can_lehmann_fsm/_0744_
+ VGND heichips25_can_lehmann_fsm/net1082 heichips25_can_lehmann_fsm/net382 sg13g2_o21ai_1
XFILLER_11_229 VPWR VGND sg13g2_decap_4
Xclkload5 clknet_leaf_3_clk clkload5/Y VPWR VGND sg13g2_inv_4
Xheichips25_can_lehmann_fsm__2487_ VGND VPWR heichips25_can_lehmann_fsm/_0926_ heichips25_can_lehmann_fsm/net395
+ heichips25_can_lehmann_fsm/_0143_ heichips25_can_lehmann_fsm/_0709_ sg13g2_a21oi_1
XFILLER_1_7 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__3039_ net774 VGND VPWR heichips25_can_lehmann_fsm/net843
+ heichips25_can_lehmann_fsm__3039_/Q clknet_leaf_19_clk sg13g2_dfrbpq_1
Xheichips25_sap3__2370_ heichips25_sap3/_1790_ VPWR heichips25_sap3/_1791_ VGND heichips25_sap3/net274
+ heichips25_sap3/net155 sg13g2_o21ai_1
XFILLER_46_137 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__4040_ heichips25_sap3/net462 VGND VPWR heichips25_sap3/_0181_ heichips25_sap3__4040_/Q
+ clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_15_513 VPWR VGND sg13g2_decap_8
XFILLER_42_354 VPWR VGND sg13g2_fill_1
XFILLER_42_343 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm_hold940 heichips25_can_lehmann_fsm__2855_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net939 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold962 heichips25_can_lehmann_fsm/_0252_ VPWR VGND heichips25_can_lehmann_fsm/net961
+ sg13g2_dlygate4sd3_1
XFILLER_24_94 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm_hold951 heichips25_can_lehmann_fsm__2932_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net950 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold984 heichips25_can_lehmann_fsm__2862_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net983 sg13g2_dlygate4sd3_1
XFILLER_10_262 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm_hold995 heichips25_can_lehmann_fsm/_0258_ VPWR VGND heichips25_can_lehmann_fsm/net994
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold973 heichips25_can_lehmann_fsm__2972_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net972 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__3001__586 VPWR VGND net585 sg13g2_tiehi
Xheichips25_sap3__3824_ heichips25_sap3/_1330_ heichips25_sap3/_1281_ heichips25_sap3__4017_/Q
+ heichips25_sap3/_1272_ heichips25_sap3__3977_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_6_255 VPWR VGND sg13g2_fill_2
XFILLER_40_82 VPWR VGND sg13g2_decap_4
XFILLER_6_288 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3755_ VPWR heichips25_sap3/_1267_ heichips25_sap3/net292 VGND sg13g2_inv_1
XFILLER_2_450 VPWR VGND sg13g2_decap_8
XFILLER_3_984 VPWR VGND sg13g2_decap_8
XFILLER_2_461 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2706_ heichips25_sap3/_0352_ heichips25_sap3/net278 heichips25_sap3__3920_/Q
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__3686_ heichips25_sap3__4005_/Q heichips25_sap3/_1066_ heichips25_sap3/net147
+ heichips25_sap3/_0146_ VPWR VGND sg13g2_mux2_1
XFILLER_49_91 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2637_ heichips25_sap3/_0300_ heichips25_sap3/_0302_ heichips25_sap3/_0303_
+ heichips25_sap3/_0304_ VPWR VGND sg13g2_nor3_1
XFILLER_2_494 VPWR VGND sg13g2_fill_1
XFILLER_27_6 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2568_ VPWR uio_out_sap3\[3\] heichips25_sap3/net45 VGND sg13g2_inv_1
X_23_ net508 uio_oe_sap3\[1\] net505 net20 VPWR VGND sg13g2_mux2_1
XFILLER_34_811 VPWR VGND sg13g2_fill_1
XFILLER_34_800 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2499_ heichips25_sap3/_1911_ VPWR heichips25_sap3/_1912_ VGND heichips25_sap3/net286
+ heichips25_sap3/net156 sg13g2_o21ai_1
XFILLER_19_874 VPWR VGND sg13g2_fill_2
XFILLER_46_682 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2410_ heichips25_can_lehmann_fsm/net491 VPWR heichips25_can_lehmann_fsm/_0671_
+ VGND heichips25_can_lehmann_fsm__2880_/Q heichips25_can_lehmann_fsm/net421 sg13g2_o21ai_1
XFILLER_21_549 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2341_ VGND VPWR heichips25_can_lehmann_fsm/_0966_ heichips25_can_lehmann_fsm/net367
+ heichips25_can_lehmann_fsm/_0070_ heichips25_can_lehmann_fsm/_0636_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2272_ VGND VPWR heichips25_can_lehmann_fsm/_1047_ heichips25_can_lehmann_fsm/_0587_
+ heichips25_can_lehmann_fsm/_0588_ heichips25_can_lehmann_fsm/net172 sg13g2_a21oi_1
XFILLER_29_17 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3873__818 VPWR net817 clkload23/A VGND sg13g2_inv_1
XFILLER_29_605 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1987_ heichips25_can_lehmann_fsm/net323 VPWR heichips25_can_lehmann_fsm/_0345_
+ VGND heichips25_can_lehmann_fsm/net1248 heichips25_can_lehmann_fsm/net177 sg13g2_o21ai_1
XFILLER_36_192 VPWR VGND sg13g2_fill_2
XFILLER_12_527 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2608_ heichips25_can_lehmann_fsm/net499 VPWR heichips25_can_lehmann_fsm/_0770_
+ VGND heichips25_can_lehmann_fsm/net897 heichips25_can_lehmann_fsm/net381 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2539_ VGND VPWR heichips25_can_lehmann_fsm/_0913_ heichips25_can_lehmann_fsm/net393
+ heichips25_can_lehmann_fsm/_0169_ heichips25_can_lehmann_fsm/_0735_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2820__567 VPWR VGND net566 sg13g2_tiehi
XFILLER_4_737 VPWR VGND sg13g2_fill_1
Xclkbuf_4_6_0_heichips25_sap3\_sap_3_inst.alu_inst.clk clknet_0_heichips25_sap3\/sap_3_inst.alu_inst.clk
+ clknet_4_6_0_heichips25_sap3\/sap_3_inst.alu_inst.clk VPWR VGND sg13g2_buf_8
XFILLER_3_269 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3540_ VGND VPWR heichips25_sap3/net96 heichips25_sap3/_1037_ heichips25_sap3/_1130_
+ heichips25_sap3/_1128_ sg13g2_a21oi_1
Xheichips25_sap3__3471_ heichips25_sap3/net57 heichips25_sap3/_1070_ heichips25_sap3/_1071_
+ heichips25_sap3/_1072_ VPWR VGND sg13g2_nor3_1
XFILLER_0_943 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2422_ heichips25_sap3/_1837_ heichips25_sap3/_1838_ heichips25_sap3/_1839_
+ VPWR VGND sg13g2_and2_1
Xheichips25_sap3__2353_ heichips25_sap3/_1774_ heichips25_sap3/_1605_ heichips25_sap3/_1515_
+ heichips25_sap3/_1549_ heichips25_sap3/net242 VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2284_ heichips25_sap3/_1701_ heichips25_sap3/_1703_ heichips25_sap3/_1704_
+ heichips25_sap3/_1705_ VPWR VGND sg13g2_nor3_1
Xheichips25_sap3__4023_ heichips25_sap3/net457 VGND VPWR heichips25_sap3/_0164_ heichips25_sap3__4023_/Q
+ clkload29/A sg13g2_dfrbpq_1
XFILLER_15_321 VPWR VGND sg13g2_decap_8
XFILLER_27_192 VPWR VGND sg13g2_decap_8
XFILLER_35_82 VPWR VGND sg13g2_fill_1
XFILLER_30_357 VPWR VGND sg13g2_fill_1
XFILLER_7_586 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__1999_ VPWR heichips25_sap3/_1425_ heichips25_sap3__3954_/Q VGND
+ sg13g2_inv_1
Xheichips25_sap3__3807_ heichips25_sap3/_1315_ heichips25_sap3/_1274_ heichips25_sap3__3943_/Q
+ heichips25_sap3/_1272_ heichips25_sap3__3975_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3738_ VGND VPWR heichips25_sap3/_1429_ heichips25_sap3/net339 heichips25_sap3/_0169_
+ heichips25_sap3/net832 sg13g2_a21oi_1
XFILLER_2_291 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3669_ heichips25_sap3/_1213_ heichips25_sap3/_0969_ heichips25_sap3/_0991_
+ VPWR VGND sg13g2_xnor2_1
Xheichips25_can_lehmann_fsm__1910_ heichips25_can_lehmann_fsm/_1216_ heichips25_can_lehmann_fsm/_1222_
+ heichips25_can_lehmann_fsm/_1162_ heichips25_can_lehmann_fsm/_1223_ VPWR VGND sg13g2_nand3_1
XFILLER_39_969 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2890_ net715 VGND VPWR heichips25_can_lehmann_fsm/_0115_
+ heichips25_can_lehmann_fsm__2890_/Q clknet_leaf_14_clk sg13g2_dfrbpq_1
XFILLER_18_2 VPWR VGND sg13g2_fill_1
X_06_ uo_out_fsm\[0\] uo_out_sap3\[0\] net507 net35 VPWR VGND sg13g2_mux2_1
Xheichips25_can_lehmann_fsm__1841_ heichips25_can_lehmann_fsm/_1155_ heichips25_can_lehmann_fsm/_1156_
+ heichips25_can_lehmann_fsm/_1154_ heichips25_can_lehmann_fsm/_1157_ VPWR VGND sg13g2_nand3_1
XFILLER_47_980 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1772_ VGND VPWR heichips25_can_lehmann_fsm__2894_/Q heichips25_can_lehmann_fsm/net296
+ heichips25_can_lehmann_fsm/_1088_ heichips25_can_lehmann_fsm/net300 sg13g2_a21oi_1
XFILLER_25_118 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm_hold1108 heichips25_can_lehmann_fsm/_0160_ VPWR VGND heichips25_can_lehmann_fsm/net1107
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1119 heichips25_can_lehmann_fsm/_0275_ VPWR VGND heichips25_can_lehmann_fsm/net1118
+ sg13g2_dlygate4sd3_1
XFILLER_33_162 VPWR VGND sg13g2_fill_1
XFILLER_21_335 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__3021__715 VPWR VGND net714 sg13g2_tiehi
Xheichips25_sap3_hold839 heichips25_sap3__4071_/A VPWR VGND heichips25_sap3/net838
+ sg13g2_dlygate4sd3_1
XFILLER_21_357 VPWR VGND sg13g2_fill_2
XFILLER_21_368 VPWR VGND sg13g2_decap_8
XFILLER_21_379 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2324_ heichips25_can_lehmann_fsm/net471 VPWR heichips25_can_lehmann_fsm/_0628_
+ VGND heichips25_can_lehmann_fsm__2836_/Q heichips25_can_lehmann_fsm/net363 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2255_ heichips25_can_lehmann_fsm/_1044_ heichips25_can_lehmann_fsm__2822_/Q
+ heichips25_can_lehmann_fsm/_0574_ VPWR VGND sg13g2_xor2_1
Xheichips25_sap3_fanout49 heichips25_sap3/_0871_ heichips25_sap3/net49 VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm__2186_ heichips25_can_lehmann_fsm/_0520_ heichips25_can_lehmann_fsm/_0519_
+ heichips25_can_lehmann_fsm/_1099_ VPWR VGND sg13g2_nand2b_1
Xoutput29 net29 uio_out[2] VPWR VGND sg13g2_buf_1
XFILLER_0_206 VPWR VGND sg13g2_decap_8
XFILLER_0_239 VPWR VGND sg13g2_decap_8
XFILLER_5_1003 VPWR VGND sg13g2_decap_8
Xheichips25_sap3_hold1163 heichips25_sap3__4030_/Q VPWR VGND heichips25_sap3/net1162
+ sg13g2_dlygate4sd3_1
XFILLER_12_324 VPWR VGND sg13g2_decap_8
XFILLER_12_346 VPWR VGND sg13g2_fill_1
XFILLER_40_699 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2976__721 VPWR VGND net720 sg13g2_tiehi
Xheichips25_sap3__2971_ heichips25_sap3/_0608_ heichips25_sap3__3907_/Q heichips25_sap3/_0607_
+ VPWR VGND sg13g2_nand2_1
XFILLER_4_523 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2872__752 VPWR VGND net751 sg13g2_tiehi
Xheichips25_sap3__3523_ heichips25_sap3/_1110_ heichips25_sap3/_1115_ heichips25_sap3/_0092_
+ VPWR VGND sg13g2_nor2b_1
XFILLER_48_733 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3454_ heichips25_sap3/_1059_ heichips25_sap3/_1056_ heichips25_sap3/_1058_
+ heichips25_sap3/net58 heichips25_sap3__3939_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3385_ heichips25_sap3/_0991_ heichips25_sap3/net59 heichips25_sap3/_0993_
+ VPWR VGND heichips25_sap3/_0969_ sg13g2_nand3b_1
Xheichips25_sap3__2405_ heichips25_sap3/_1813_ heichips25_sap3/_1816_ heichips25_sap3/_1823_
+ uio_out_sap3\[6\] VPWR VGND heichips25_sap3/_1812_ sg13g2_nand4_1
Xheichips25_sap3__2336_ heichips25_sap3/_1486_ VPWR heichips25_sap3/_1757_ VGND heichips25_sap3/_1363_
+ heichips25_sap3/_1553_ sg13g2_o21ai_1
XFILLER_46_81 VPWR VGND sg13g2_fill_1
XFILLER_16_630 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2267_ heichips25_sap3/_1688_ heichips25_sap3/_1441_ heichips25_sap3/_1662_
+ VPWR VGND sg13g2_nand2_1
XFILLER_15_151 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2198_ heichips25_sap3/_1434_ heichips25_sap3/net268 heichips25_sap3/_1619_
+ VPWR VGND heichips25_sap3/net270 sg13g2_nand3b_1
XFILLER_15_184 VPWR VGND sg13g2_decap_8
XFILLER_15_195 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__4006_ heichips25_sap3/net443 VGND VPWR heichips25_sap3/_0147_ heichips25_sap3__4006_/Q
+ heichips25_sap3__4009_/CLK sg13g2_dfrbpq_1
XFILLER_30_176 VPWR VGND sg13g2_decap_8
XFILLER_30_187 VPWR VGND sg13g2_fill_2
XFILLER_7_42 VPWR VGND sg13g2_fill_2
XFILLER_11_390 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2955__805 VPWR VGND net804 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2040_ VGND VPWR heichips25_can_lehmann_fsm/net177 heichips25_can_lehmann_fsm/_0388_
+ heichips25_can_lehmann_fsm/_0016_ heichips25_can_lehmann_fsm/_0389_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2918__660 VPWR VGND net659 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2942_ net567 VGND VPWR heichips25_can_lehmann_fsm/net971
+ heichips25_can_lehmann_fsm__2942_/Q clknet_leaf_19_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2873_ net749 VGND VPWR heichips25_can_lehmann_fsm/net1067
+ heichips25_can_lehmann_fsm__2873_/Q clknet_leaf_0_clk sg13g2_dfrbpq_1
XFILLER_27_917 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1824_ heichips25_can_lehmann_fsm__3045_/Q heichips25_can_lehmann_fsm__3044_/Q
+ heichips25_can_lehmann_fsm/_1140_ VPWR VGND sg13g2_nor2_1
Xclkbuf_leaf_18_clk clknet_2_2__leaf_clk clknet_leaf_18_clk VPWR VGND sg13g2_buf_8
Xheichips25_can_lehmann_fsm__2849__798 VPWR VGND net797 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__1755_ heichips25_can_lehmann_fsm/_0979_ heichips25_can_lehmann_fsm/_0980_
+ heichips25_can_lehmann_fsm/_0978_ heichips25_can_lehmann_fsm/_1075_ VPWR VGND heichips25_can_lehmann_fsm/_1071_
+ sg13g2_nand4_1
Xheichips25_can_lehmann_fsm__1686_ heichips25_can_lehmann_fsm/_1009_ VPWR heichips25_can_lehmann_fsm/_1010_
+ VGND heichips25_can_lehmann_fsm__2873_/Q heichips25_can_lehmann_fsm/net336 sg13g2_o21ai_1
XFILLER_21_121 VPWR VGND sg13g2_fill_1
XFILLER_34_471 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2307_ heichips25_can_lehmann_fsm/_0616_ heichips25_can_lehmann_fsm__2832_/Q
+ heichips25_can_lehmann_fsm/_1052_ VPWR VGND sg13g2_xnor2_1
Xheichips25_can_lehmann_fsm__2238_ VGND VPWR heichips25_can_lehmann_fsm/net205 heichips25_can_lehmann_fsm/_0559_
+ heichips25_can_lehmann_fsm/_0043_ heichips25_can_lehmann_fsm/_0560_ sg13g2_a21oi_1
Xheichips25_sap3__3879__824 VPWR net823 heichips25_sap3__3996_/CLK VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__2169_ heichips25_can_lehmann_fsm/net1215 VPWR heichips25_can_lehmann_fsm/_0506_
+ VGND heichips25_can_lehmann_fsm__2803_/Q heichips25_can_lehmann_fsm__2802_/Q sg13g2_o21ai_1
XFILLER_29_276 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3170_ heichips25_sap3/_0783_ heichips25_sap3/net104 heichips25_sap3__3954_/Q
+ heichips25_sap3/net109 heichips25_sap3__3962_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2121_ heichips25_sap3__3928_/Q heichips25_sap3__3892_/Q heichips25_sap3__3890_/Q
+ heichips25_sap3/net254 heichips25_sap3__3891_/Q heichips25_sap3/net263 heichips25_sap3/_1542_
+ VPWR VGND sg13g2_mux4_1
XFILLER_25_460 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2052_ heichips25_sap3/_1472_ heichips25_sap3/net237 heichips25_sap3/net248
+ heichips25_sap3/_1473_ VPWR VGND sg13g2_a21o_1
XFILLER_12_176 VPWR VGND sg13g2_decap_4
XFILLER_8_158 VPWR VGND sg13g2_decap_4
XFILLER_32_72 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2954_ heichips25_sap3/_0592_ heichips25_sap3/_1374_ heichips25_sap3/_0442_
+ VPWR VGND sg13g2_nand2_1
XFILLER_5_887 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2885_ heichips25_sap3/_0525_ VPWR heichips25_sap3/_0526_ VGND heichips25_sap3/net280
+ heichips25_sap3/_0441_ sg13g2_o21ai_1
Xheichips25_sap3__3506_ heichips25_sap3/_1101_ net44 heichips25_sap3/_1088_ VPWR VGND
+ sg13g2_nand2_1
Xheichips25_sap3__3437_ heichips25_sap3/_0999_ heichips25_sap3/_1015_ heichips25_sap3/_1043_
+ VPWR VGND heichips25_sap3/_1036_ sg13g2_nand3b_1
Xheichips25_sap3__3368_ heichips25_sap3/_0977_ heichips25_sap3/_0952_ heichips25_sap3/_0966_
+ VPWR VGND sg13g2_xnor2_1
X_15__517 VPWR VGND net516 sg13g2_tielo
XFILLER_16_460 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2319_ heichips25_sap3/_1740_ heichips25_sap3/_1680_ heichips25_sap3/_1713_
+ heichips25_sap3/_1732_ VPWR VGND sg13g2_and3_1
Xheichips25_sap3__3299_ heichips25_sap3/_0909_ heichips25_sap3/_0910_ heichips25_sap3/_0911_
+ VPWR VGND sg13g2_and2_1
Xheichips25_can_lehmann_fsm__1540_ VPWR heichips25_can_lehmann_fsm/_0864_ heichips25_can_lehmann_fsm/net1164
+ VGND sg13g2_inv_1
XFILLER_32_920 VPWR VGND sg13g2_fill_1
XFILLER_32_975 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_7_clk clknet_2_1__leaf_clk clknet_leaf_7_clk VPWR VGND sg13g2_buf_8
Xheichips25_can_lehmann_fsm__2023_ VGND VPWR heichips25_can_lehmann_fsm/net1244 heichips25_can_lehmann_fsm/net188
+ heichips25_can_lehmann_fsm/_0375_ heichips25_can_lehmann_fsm/net191 sg13g2_a21oi_1
XFILLER_37_28 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2925_ net635 VGND VPWR heichips25_can_lehmann_fsm/_0150_
+ heichips25_can_lehmann_fsm__2925_/Q clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_2_1028 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2856_ net783 VGND VPWR heichips25_can_lehmann_fsm/_0081_
+ heichips25_can_lehmann_fsm__2856_/Q clknet_leaf_10_clk sg13g2_dfrbpq_1
XFILLER_26_224 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1807_ heichips25_can_lehmann_fsm/_1114_ heichips25_can_lehmann_fsm/_1122_
+ heichips25_can_lehmann_fsm/_1123_ VPWR VGND sg13g2_nor2_1
Xheichips25_can_lehmann_fsm__2787_ net632 VGND VPWR heichips25_can_lehmann_fsm/net1241
+ heichips25_can_lehmann_fsm__2787_/Q clknet_leaf_1_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1738_ VGND VPWR heichips25_can_lehmann_fsm/_1058_ heichips25_can_lehmann_fsm/_1057_
+ heichips25_can_lehmann_fsm/_1056_ sg13g2_or2_1
Xheichips25_can_lehmann_fsm__1669_ heichips25_can_lehmann_fsm/net338 heichips25_can_lehmann_fsm/_0992_
+ heichips25_can_lehmann_fsm/_0993_ VPWR VGND sg13g2_and2_1
Xheichips25_sap3__2670_ VPWR VGND heichips25_sap3/_1848_ heichips25_sap3/net66 heichips25_sap3/_1851_
+ heichips25_sap3/_1400_ uio_oe_sap3\[4\] heichips25_sap3/net90 sg13g2_a221oi_1
XFILLER_2_857 VPWR VGND sg13g2_fill_1
XFILLER_2_868 VPWR VGND sg13g2_fill_2
XFILLER_1_345 VPWR VGND sg13g2_fill_1
XFILLER_49_338 VPWR VGND sg13g2_fill_1
XFILLER_45_544 VPWR VGND sg13g2_decap_8
XFILLER_45_533 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3222_ heichips25_sap3/_0831_ heichips25_sap3/_0832_ heichips25_sap3/_0833_
+ heichips25_sap3/_0834_ heichips25_sap3/_0835_ VPWR VGND sg13g2_and4_1
XFILLER_45_577 VPWR VGND sg13g2_fill_1
XFILLER_17_279 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3153_ heichips25_sap3/_0667_ heichips25_sap3/_0679_ heichips25_sap3/_0697_
+ heichips25_sap3/_0766_ VPWR VGND sg13g2_nor3_1
XFILLER_32_205 VPWR VGND sg13g2_fill_1
Xclkbuf_5_9__f_heichips25_sap3\_sap_3_inst.alu_inst.clk heichips25_sap3__4018_/CLK
+ clknet_4_4_0_heichips25_sap3\/sap_3_inst.alu_inst.clk VPWR VGND sg13g2_buf_16
Xheichips25_sap3__2104_ heichips25_sap3/_1514_ heichips25_sap3/_1519_ heichips25_sap3/_1504_
+ heichips25_sap3/_1525_ VPWR VGND heichips25_sap3/_1523_ sg13g2_nand4_1
XFILLER_41_761 VPWR VGND sg13g2_fill_1
XFILLER_14_964 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3084_ heichips25_sap3/_0690_ heichips25_sap3/_0695_ heichips25_sap3/_1753_
+ heichips25_sap3/_0697_ VPWR VGND sg13g2_nand3_1
Xheichips25_sap3__2035_ VPWR heichips25_sap3/_1456_ heichips25_sap3/_1455_ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__3004__562 VPWR VGND net561 sg13g2_tiehi
Xheichips25_can_lehmann_fsm_hold1280 heichips25_can_lehmann_fsm__2814_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1279 sg13g2_dlygate4sd3_1
XFILLER_9_478 VPWR VGND sg13g2_decap_4
XFILLER_9_489 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3986_ heichips25_sap3/net441 VGND VPWR heichips25_sap3/_0127_ heichips25_sap3__3986_/Q
+ clkload20/A sg13g2_dfrbpq_1
Xheichips25_sap3__2937_ heichips25_sap3/_0576_ heichips25_sap3/net276 heichips25_sap3/net211
+ VPWR VGND sg13g2_xnor2_1
Xheichips25_sap3__2868_ heichips25_sap3/_0510_ heichips25_sap3/_0417_ heichips25_sap3/net285
+ heichips25_sap3/_0359_ heichips25_sap3/net159 VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2799_ heichips25_sap3/_0344_ heichips25_sap3/_0443_ heichips25_sap3/_0444_
+ VPWR VGND sg13g2_and2_1
XFILLER_49_872 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2710_ heichips25_can_lehmann_fsm/net486 VPWR heichips25_can_lehmann_fsm/_0821_
+ VGND heichips25_can_lehmann_fsm/net1029 heichips25_can_lehmann_fsm/net378 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2641_ VGND VPWR heichips25_can_lehmann_fsm/_0887_ heichips25_can_lehmann_fsm/net360
+ heichips25_can_lehmann_fsm/_0220_ heichips25_can_lehmann_fsm/_0786_ sg13g2_a21oi_1
XFILLER_24_706 VPWR VGND sg13g2_fill_2
XFILLER_36_599 VPWR VGND sg13g2_decap_8
XFILLER_17_780 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2572_ heichips25_can_lehmann_fsm/net482 VPWR heichips25_can_lehmann_fsm/_0752_
+ VGND heichips25_can_lehmann_fsm__2960_/Q heichips25_can_lehmann_fsm/net374 sg13g2_o21ai_1
XFILLER_23_19 VPWR VGND sg13g2_fill_2
XFILLER_31_271 VPWR VGND sg13g2_decap_8
XFILLER_31_282 VPWR VGND sg13g2_fill_2
XFILLER_2_109 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__3055_ net670 VGND VPWR heichips25_can_lehmann_fsm/net1044
+ heichips25_can_lehmann_fsm__3055_/Q clknet_leaf_15_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2006_ heichips25_can_lehmann_fsm/net321 VPWR heichips25_can_lehmann_fsm/_0361_
+ VGND heichips25_can_lehmann_fsm__2786_/Q heichips25_can_lehmann_fsm/net178 sg13g2_o21ai_1
XFILLER_24_1007 VPWR VGND sg13g2_fill_1
XFILLER_46_308 VPWR VGND sg13g2_decap_8
XFILLER_39_360 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2908_ net679 VGND VPWR heichips25_can_lehmann_fsm/_0133_
+ heichips25_can_lehmann_fsm__2908_/Q clknet_leaf_12_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2839_ net528 VGND VPWR heichips25_can_lehmann_fsm/_0064_
+ heichips25_can_lehmann_fsm__2839_/Q clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_14_238 VPWR VGND sg13g2_fill_1
XFILLER_15_739 VPWR VGND sg13g2_fill_2
XFILLER_7_938 VPWR VGND sg13g2_decap_4
XFILLER_6_426 VPWR VGND sg13g2_decap_8
XFILLER_13_63 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3840_ heichips25_sap3/_0181_ heichips25_sap3/net1197 heichips25_sap3/_0018_
+ VPWR VGND sg13g2_xnor2_1
XFILLER_6_437 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3771_ heichips25_sap3/_1283_ heichips25_sap3/_1282_ heichips25_sap3__3947_/Q
+ heichips25_sap3/_1281_ heichips25_sap3__4011_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2722_ VGND VPWR heichips25_sap3/_0356_ heichips25_sap3/_0367_ heichips25_sap3/_0368_
+ heichips25_sap3/_0354_ sg13g2_a21oi_1
XFILLER_2_643 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__3034__566 VPWR VGND net565 sg13g2_tiehi
XFILLER_49_102 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2653_ heichips25_sap3/net249 heichips25_sap3/net248 heichips25_sap3/_0319_
+ heichips25_sap3/_0320_ VPWR VGND sg13g2_nor3_1
XFILLER_1_153 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2584_ heichips25_sap3/_1654_ heichips25_sap3/_0247_ heichips25_sap3/_0256_
+ heichips25_sap3/_0257_ VPWR VGND sg13g2_nor3_1
Xheichips25_can_lehmann_fsm__2830__547 VPWR VGND net546 sg13g2_tiehi
XFILLER_38_93 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3205_ heichips25_sap3/_0818_ heichips25_sap3__3942_/Q heichips25_sap3/net128
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__3136_ heichips25_sap3/_0731_ heichips25_sap3/net166 heichips25_sap3/_0749_
+ VPWR VGND sg13g2_and2_1
Xheichips25_sap3__3067_ heichips25_sap3/_0666_ heichips25_sap3/_0679_ heichips25_sap3/_0680_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__2018_ VGND VPWR heichips25_sap3/_1439_ heichips25_sap3/net269 heichips25_sap3/net272
+ sg13g2_or2_1
XFILLER_9_220 VPWR VGND sg13g2_decap_8
XFILLER_9_231 VPWR VGND sg13g2_fill_1
Xclkload23 VPWR clkload23/Y clkload23/A VGND sg13g2_inv_1
Xclkload12 VPWR clkload12/Y clknet_leaf_20_clk VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm_fanout329 heichips25_can_lehmann_fsm/net330 heichips25_can_lehmann_fsm/net329
+ VPWR VGND sg13g2_buf_1
Xheichips25_sap3__3969_ heichips25_sap3/net440 VGND VPWR heichips25_sap3/_0110_ heichips25_sap3__3969_/Q
+ heichips25_sap3__4017_/CLK sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm_fanout318 heichips25_can_lehmann_fsm/net320 heichips25_can_lehmann_fsm/net318
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout307 heichips25_can_lehmann_fsm/net309 heichips25_can_lehmann_fsm/net307
+ VPWR VGND sg13g2_buf_1
XFILLER_36_385 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2624_ heichips25_can_lehmann_fsm/net482 VPWR heichips25_can_lehmann_fsm/_0778_
+ VGND heichips25_can_lehmann_fsm__2986_/Q heichips25_can_lehmann_fsm/net374 sg13g2_o21ai_1
XFILLER_24_569 VPWR VGND sg13g2_fill_1
XFILLER_34_29 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2555_ VGND VPWR heichips25_can_lehmann_fsm/_0909_ heichips25_can_lehmann_fsm/net407
+ heichips25_can_lehmann_fsm/_0177_ heichips25_can_lehmann_fsm/_0743_ sg13g2_a21oi_1
Xclkload6 VPWR clkload6/Y clknet_leaf_4_clk VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__2486_ heichips25_can_lehmann_fsm/net476 VPWR heichips25_can_lehmann_fsm/_0709_
+ VGND heichips25_can_lehmann_fsm/net1070 heichips25_can_lehmann_fsm/net395 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__3038_ net790 VGND VPWR heichips25_can_lehmann_fsm/_0263_
+ heichips25_can_lehmann_fsm__3038_/Q clknet_leaf_19_clk sg13g2_dfrbpq_1
XFILLER_15_503 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__3029__646 VPWR VGND net645 sg13g2_tiehi
XFILLER_27_341 VPWR VGND sg13g2_fill_1
XFILLER_28_886 VPWR VGND sg13g2_decap_8
XFILLER_42_311 VPWR VGND sg13g2_decap_8
XFILLER_15_569 VPWR VGND sg13g2_decap_8
XFILLER_24_51 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm_hold941 heichips25_can_lehmann_fsm/_0080_ VPWR VGND heichips25_can_lehmann_fsm/net940
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold930 heichips25_can_lehmann_fsm/_0220_ VPWR VGND heichips25_can_lehmann_fsm/net929
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold952 heichips25_can_lehmann_fsm__3030_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net951 sg13g2_dlygate4sd3_1
XFILLER_10_230 VPWR VGND sg13g2_decap_8
XFILLER_10_241 VPWR VGND sg13g2_fill_2
XFILLER_11_753 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm_hold963 heichips25_can_lehmann_fsm__2922_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net962 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold974 heichips25_can_lehmann_fsm__2890_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net973 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold985 heichips25_can_lehmann_fsm__2984_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net984 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold996 heichips25_can_lehmann_fsm__2993_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net995 sg13g2_dlygate4sd3_1
Xheichips25_sap3__3823_ heichips25_sap3/_1329_ heichips25_sap3/_1279_ heichips25_sap3__3969_/Q
+ heichips25_sap3/_1274_ heichips25_sap3__3945_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_40_94 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3754_ heichips25_sap3__4043_/Q heichips25_sap3__4042_/Q heichips25_sap3/_1260_
+ heichips25_sap3/_1266_ VPWR VGND sg13g2_nor3_1
XFILLER_3_963 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2705_ heichips25_sap3/net278 heichips25_sap3__3920_/Q heichips25_sap3/_0351_
+ VPWR VGND sg13g2_and2_1
Xheichips25_sap3__3685_ heichips25_sap3__4004_/Q heichips25_sap3/_1175_ heichips25_sap3/net147
+ heichips25_sap3/_0145_ VPWR VGND sg13g2_mux2_1
Xheichips25_sap3__2636_ heichips25_sap3/_1725_ heichips25_sap3/_0296_ heichips25_sap3/_1621_
+ heichips25_sap3/_0303_ VPWR VGND heichips25_sap3/_0298_ sg13g2_nand4_1
X_22_ net uio_oe_sap3\[0\] net505 net19 VPWR VGND sg13g2_mux2_1
XFILLER_1_33 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2567_ heichips25_sap3/_0232_ heichips25_sap3/_0234_ heichips25_sap3/_0241_
+ heichips25_sap3/_0242_ VPWR VGND sg13g2_nor3_1
XFILLER_46_661 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2498_ heichips25_sap3/_1911_ heichips25_sap3/net156 heichips25_sap3/_1910_
+ VPWR VGND sg13g2_nand2_1
XFILLER_18_341 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2882__732 VPWR VGND net731 sg13g2_tiehi
XFILLER_21_528 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3119_ VPWR heichips25_sap3/_0732_ heichips25_sap3/_0731_ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__2340_ heichips25_can_lehmann_fsm/net474 VPWR heichips25_can_lehmann_fsm/_0636_
+ VGND heichips25_can_lehmann_fsm__2844_/Q heichips25_can_lehmann_fsm/net367 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2271_ heichips25_can_lehmann_fsm/_0587_ heichips25_can_lehmann_fsm/net1182
+ heichips25_can_lehmann_fsm/_1046_ VPWR VGND sg13g2_nand2b_1
Xclkbuf_5_27__f_heichips25_sap3\_sap_3_inst.alu_inst.clk clkload27/A clknet_4_13_0_heichips25_sap3\/sap_3_inst.alu_inst.clk
+ VPWR VGND sg13g2_buf_16
Xheichips25_can_lehmann_fsm__1986_ heichips25_can_lehmann_fsm/_0343_ heichips25_can_lehmann_fsm/_0341_
+ heichips25_can_lehmann_fsm/_0342_ heichips25_can_lehmann_fsm/_0344_ VPWR VGND sg13g2_a21o_1
XFILLER_36_171 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2783__641 VPWR VGND net640 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2607_ VGND VPWR heichips25_can_lehmann_fsm/_0896_ heichips25_can_lehmann_fsm/net422
+ heichips25_can_lehmann_fsm/_0203_ heichips25_can_lehmann_fsm/_0769_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2538_ heichips25_can_lehmann_fsm/net466 VPWR heichips25_can_lehmann_fsm/_0735_
+ VGND heichips25_can_lehmann_fsm/net969 heichips25_can_lehmann_fsm/net393 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2469_ VGND VPWR heichips25_can_lehmann_fsm/_0930_ heichips25_can_lehmann_fsm/net377
+ heichips25_can_lehmann_fsm/_0134_ heichips25_can_lehmann_fsm/_0700_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2859__778 VPWR VGND net777 sg13g2_tiehi
XFILLER_0_922 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3470_ VGND VPWR heichips25_sap3/_0764_ heichips25_sap3/_0973_ heichips25_sap3/_1071_
+ heichips25_sap3/_0863_ sg13g2_a21oi_1
Xheichips25_sap3__2421_ heichips25_sap3/_1838_ heichips25_sap3/net72 heichips25_sap3__3984_/Q
+ heichips25_sap3/_1744_ heichips25_sap3__3992_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_0_999 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2352_ heichips25_sap3/_1480_ heichips25_sap3/_1619_ heichips25_sap3/_1773_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__2283_ heichips25_sap3/_1364_ heichips25_sap3/_1621_ heichips25_sap3/_1645_
+ heichips25_sap3/_1704_ VPWR VGND sg13g2_nor3_1
XFILLER_27_160 VPWR VGND sg13g2_decap_8
XFILLER_27_171 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__4022_ heichips25_sap3/net457 VGND VPWR heichips25_sap3/_0163_ heichips25_sap3__4022_/Q
+ clkload28/A sg13g2_dfrbpq_1
XFILLER_37_1028 VPWR VGND sg13g2_fill_1
XFILLER_42_196 VPWR VGND sg13g2_decap_8
XFILLER_7_521 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__1998_ VPWR heichips25_sap3/_1424_ heichips25_sap3__3970_/Q VGND
+ sg13g2_inv_1
Xheichips25_sap3__3806_ heichips25_sap3/_1314_ heichips25_sap3/_1279_ heichips25_sap3__3967_/Q
+ heichips25_sap3/net292 heichips25_sap3__3959_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3737_ VGND VPWR heichips25_sap3/_1246_ heichips25_sap3/_1253_ heichips25_sap3/_0168_
+ heichips25_sap3/_1247_ sg13g2_a21oi_1
Xheichips25_sap3__3668_ heichips25_sap3/net828 heichips25_sap3/net111 heichips25_sap3/_1212_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__2619_ heichips25_sap3/_0001_ heichips25_sap3/_1366_ heichips25_sap3/_0288_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__3599_ VGND VPWR heichips25_sap3/net60 heichips25_sap3/net99 heichips25_sap3/_1172_
+ heichips25_sap3/net94 sg13g2_a21oi_1
X_05_ net2 net1 _01_ VPWR VGND sg13g2_and2_1
Xheichips25_can_lehmann_fsm__1840_ heichips25_can_lehmann_fsm/_1156_ heichips25_can_lehmann_fsm__3058_/Q
+ heichips25_can_lehmann_fsm/net354 VPWR VGND sg13g2_xnor2_1
XFILLER_26_609 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1771_ heichips25_can_lehmann_fsm/_1087_ heichips25_can_lehmann_fsm/net294
+ heichips25_can_lehmann_fsm__2966_/Q heichips25_can_lehmann_fsm/net305 heichips25_can_lehmann_fsm__2942_/Q
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2947__548 VPWR VGND net547 sg13g2_tiehi
XFILLER_18_182 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_hold1109 heichips25_can_lehmann_fsm__2917_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1108 sg13g2_dlygate4sd3_1
XFILLER_22_859 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2323_ VGND VPWR heichips25_can_lehmann_fsm/_0971_ heichips25_can_lehmann_fsm/net403
+ heichips25_can_lehmann_fsm/_0061_ heichips25_can_lehmann_fsm/_0627_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2254_ VGND VPWR heichips25_can_lehmann_fsm/net206 heichips25_can_lehmann_fsm/_0572_
+ heichips25_can_lehmann_fsm/_0046_ heichips25_can_lehmann_fsm/_0573_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2185_ heichips25_can_lehmann_fsm/net1210 VPWR heichips25_can_lehmann_fsm/_0519_
+ VGND heichips25_can_lehmann_fsm__2806_/Q heichips25_can_lehmann_fsm/_1098_ sg13g2_o21ai_1
Xoutput19 net19 uio_oe[0] VPWR VGND sg13g2_buf_1
XFILLER_0_229 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1969_ VPWR VGND heichips25_can_lehmann_fsm/_0327_ heichips25_can_lehmann_fsm/_0328_
+ heichips25_can_lehmann_fsm/net184 heichips25_can_lehmann_fsm/net1249 heichips25_can_lehmann_fsm/_0329_
+ heichips25_can_lehmann_fsm/net197 sg13g2_a221oi_1
XFILLER_16_119 VPWR VGND sg13g2_fill_1
Xheichips25_sap3_hold1131 heichips25_sap3__4061_/Q VPWR VGND heichips25_sap3/net1130
+ sg13g2_dlygate4sd3_1
Xheichips25_sap3_hold1120 heichips25_sap3__4052_/Q VPWR VGND heichips25_sap3/net1119
+ sg13g2_dlygate4sd3_1
XFILLER_12_303 VPWR VGND sg13g2_decap_8
Xheichips25_sap3_hold1164 heichips25_sap3/_1255_ VPWR VGND heichips25_sap3/net1163
+ sg13g2_dlygate4sd3_1
XFILLER_24_174 VPWR VGND sg13g2_fill_2
Xheichips25_sap3_hold1142 heichips25_sap3__4033_/Q VPWR VGND heichips25_sap3/net1141
+ sg13g2_dlygate4sd3_1
XFILLER_8_318 VPWR VGND sg13g2_decap_8
XFILLER_8_307 VPWR VGND sg13g2_fill_2
XFILLER_12_358 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2970_ heichips25_sap3/net167 heichips25_sap3/net153 heichips25_sap3/_0607_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__3522_ heichips25_sap3/_1111_ heichips25_sap3/_1113_ heichips25_sap3/net109
+ heichips25_sap3/_1115_ VPWR VGND heichips25_sap3/_1114_ sg13g2_nand4_1
Xheichips25_can_lehmann_fsm_fanout490 heichips25_can_lehmann_fsm/net503 heichips25_can_lehmann_fsm/net490
+ VPWR VGND sg13g2_buf_1
XFILLER_47_222 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3453_ heichips25_sap3/net58 heichips25_sap3/_1057_ heichips25_sap3/_1058_
+ VPWR VGND sg13g2_nor2b_1
Xheichips25_sap3__3384_ heichips25_sap3/_0992_ heichips25_sap3/_0991_ heichips25_sap3/_0969_
+ VPWR VGND sg13g2_nand2b_1
Xheichips25_sap3__2404_ heichips25_sap3/_1822_ heichips25_sap3/_1818_ heichips25_sap3/net66
+ heichips25_sap3/_1823_ VPWR VGND sg13g2_a21o_1
XFILLER_46_60 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2335_ heichips25_sap3/_1756_ heichips25_sap3/_1755_ heichips25_sap3/_1486_
+ heichips25_sap3/_1754_ heichips25_sap3/_1685_ VPWR VGND sg13g2_a22oi_1
XFILLER_29_981 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2266_ heichips25_sap3/_1687_ heichips25_sap3/_1685_ heichips25_sap3/_1686_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__2197_ heichips25_sap3/_1362_ heichips25_sap3/net270 heichips25_sap3/_1435_
+ heichips25_sap3/_1618_ VPWR VGND sg13g2_nor3_1
Xheichips25_sap3__4005_ heichips25_sap3/net449 VGND VPWR heichips25_sap3/_0146_ heichips25_sap3__4005_/Q
+ heichips25_sap3__4005_/CLK sg13g2_dfrbpq_1
XFILLER_31_623 VPWR VGND sg13g2_fill_2
XFILLER_31_645 VPWR VGND sg13g2_fill_2
XFILLER_8_841 VPWR VGND sg13g2_decap_4
XFILLER_12_881 VPWR VGND sg13g2_fill_2
XFILLER_7_65 VPWR VGND sg13g2_decap_4
XFILLER_7_98 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2941_ net571 VGND VPWR heichips25_can_lehmann_fsm/_0166_
+ heichips25_can_lehmann_fsm__2941_/Q clknet_leaf_18_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2872_ net751 VGND VPWR heichips25_can_lehmann_fsm/_0097_
+ heichips25_can_lehmann_fsm__2872_/Q clknet_leaf_22_clk sg13g2_dfrbpq_1
XFILLER_16_0 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1823_ heichips25_can_lehmann_fsm/_1137_ heichips25_can_lehmann_fsm/_1136_
+ heichips25_can_lehmann_fsm/_1133_ heichips25_can_lehmann_fsm/_1139_ VPWR VGND sg13g2_a21o_1
Xheichips25_can_lehmann_fsm__1754_ heichips25_can_lehmann_fsm__2792_/Q heichips25_can_lehmann_fsm__2791_/Q
+ heichips25_can_lehmann_fsm__2790_/Q heichips25_can_lehmann_fsm/_1072_ heichips25_can_lehmann_fsm/_1074_
+ VPWR VGND sg13g2_nor4_1
Xheichips25_can_lehmann_fsm__1685_ heichips25_can_lehmann_fsm/_1006_ heichips25_can_lehmann_fsm/_1007_
+ heichips25_can_lehmann_fsm/_1005_ heichips25_can_lehmann_fsm/_1009_ VPWR VGND heichips25_can_lehmann_fsm/_1008_
+ sg13g2_nand4_1
XFILLER_21_155 VPWR VGND sg13g2_fill_2
XFILLER_21_188 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2306_ VGND VPWR heichips25_can_lehmann_fsm/net209 heichips25_can_lehmann_fsm/_0614_
+ heichips25_can_lehmann_fsm/_0056_ heichips25_can_lehmann_fsm/_0615_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2237_ heichips25_can_lehmann_fsm/net329 VPWR heichips25_can_lehmann_fsm/_0560_
+ VGND heichips25_can_lehmann_fsm/net1212 heichips25_can_lehmann_fsm/net205 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2168_ VGND VPWR heichips25_can_lehmann_fsm/_0503_ heichips25_can_lehmann_fsm/_0504_
+ heichips25_can_lehmann_fsm/_0028_ heichips25_can_lehmann_fsm/_0505_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2099_ heichips25_can_lehmann_fsm/net323 VPWR heichips25_can_lehmann_fsm/_0440_
+ VGND heichips25_can_lehmann_fsm/net344 heichips25_can_lehmann_fsm/net179 sg13g2_o21ai_1
Xheichips25_sap3__2120_ heichips25_sap3/_1364_ heichips25_sap3__3928_/Q heichips25_sap3/_1541_
+ VPWR VGND sg13g2_nor2_1
XFILLER_41_921 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2051_ heichips25_sap3/net257 heichips25_sap3/_1435_ heichips25_sap3/_1439_
+ heichips25_sap3/_1444_ heichips25_sap3/_1472_ VPWR VGND sg13g2_nor4_1
XFILLER_12_144 VPWR VGND sg13g2_decap_4
XFILLER_8_126 VPWR VGND sg13g2_fill_2
XFILLER_12_199 VPWR VGND sg13g2_decap_8
XFILLER_5_833 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2953_ heichips25_sap3/_1892_ heichips25_sap3/_1896_ heichips25_sap3/net254
+ heichips25_sap3/_0591_ VPWR VGND sg13g2_nand3_1
XFILLER_4_310 VPWR VGND sg13g2_fill_2
XFILLER_5_877 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2884_ heichips25_sap3/_0525_ heichips25_sap3/_0417_ heichips25_sap3/net282
+ heichips25_sap3/_0416_ heichips25_sap3/net278 VPWR VGND sg13g2_a22oi_1
XFILLER_4_387 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3505_ heichips25_sap3/_1100_ heichips25_sap3/net122 heichips25_sap3/_0923_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__3436_ heichips25_sap3/_1036_ VPWR heichips25_sap3/_1042_ VGND heichips25_sap3/_1000_
+ heichips25_sap3/_1014_ sg13g2_o21ai_1
Xheichips25_sap3__3367_ heichips25_sap3/_0857_ heichips25_sap3/_0951_ heichips25_sap3/net53
+ heichips25_sap3/_0976_ VPWR VGND heichips25_sap3/_0966_ sg13g2_nand4_1
XFILLER_35_236 VPWR VGND sg13g2_fill_1
XFILLER_35_258 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2318_ heichips25_sap3/_1680_ heichips25_sap3/_1693_ heichips25_sap3/_1713_
+ heichips25_sap3/_1732_ heichips25_sap3/_1739_ VPWR VGND sg13g2_nor4_1
Xheichips25_sap3__3298_ heichips25_sap3/net48 heichips25_sap3/net59 heichips25_sap3/net51
+ heichips25_sap3/_0910_ VPWR VGND sg13g2_a21o_1
Xheichips25_sap3__2249_ heichips25_sap3/net250 heichips25_sap3/_1460_ heichips25_sap3/_1518_
+ heichips25_sap3/_1670_ VPWR VGND sg13g2_nor3_1
Xheichips25_can_lehmann_fsm__2840__527 VPWR VGND net526 sg13g2_tiehi
XFILLER_7_170 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2022_ heichips25_can_lehmann_fsm/_0374_ heichips25_can_lehmann_fsm/_1072_
+ heichips25_can_lehmann_fsm/_0373_ VPWR VGND sg13g2_nand2_1
Xheichips25_can_lehmann_fsm__2924_ net639 VGND VPWR heichips25_can_lehmann_fsm/net894
+ heichips25_can_lehmann_fsm__2924_/Q clknet_leaf_0_clk sg13g2_dfrbpq_1
XFILLER_2_1007 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2855_ net785 VGND VPWR heichips25_can_lehmann_fsm/net940
+ heichips25_can_lehmann_fsm__2855_/Q clknet_leaf_9_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1806_ heichips25_can_lehmann_fsm/_1122_ heichips25_can_lehmann_fsm/_1116_
+ heichips25_can_lehmann_fsm/_1121_ heichips25_can_lehmann_fsm/net301 heichips25_can_lehmann_fsm/_0950_
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2786_ net634 VGND VPWR heichips25_can_lehmann_fsm/net1243
+ heichips25_can_lehmann_fsm__2786_/Q clknet_leaf_1_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1737_ VGND VPWR heichips25_can_lehmann_fsm/_1057_ heichips25_can_lehmann_fsm/net345
+ heichips25_can_lehmann_fsm__2799_/Q sg13g2_or2_1
XFILLER_23_910 VPWR VGND sg13g2_fill_1
XFILLER_23_943 VPWR VGND sg13g2_fill_1
XFILLER_22_431 VPWR VGND sg13g2_decap_4
XFILLER_10_615 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1668_ heichips25_can_lehmann_fsm/net353 heichips25_can_lehmann_fsm/net351
+ heichips25_can_lehmann_fsm/_0992_ VPWR VGND sg13g2_nor2b_1
Xheichips25_can_lehmann_fsm__1599_ VPWR heichips25_can_lehmann_fsm/_0923_ heichips25_can_lehmann_fsm/net893
+ VGND sg13g2_inv_1
XFILLER_5_129 VPWR VGND sg13g2_decap_8
XFILLER_49_317 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3221_ heichips25_sap3/_0834_ heichips25_sap3/net133 heichips25_sap3__3997_/Q
+ heichips25_sap3/net134 heichips25_sap3__3973_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_27_51 VPWR VGND sg13g2_fill_1
XFILLER_27_73 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3152_ heichips25_sap3/_0765_ heichips25_sap3__3939_/Q heichips25_sap3/net105
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__2103_ heichips25_sap3/_1504_ heichips25_sap3/_1514_ heichips25_sap3/_1519_
+ heichips25_sap3/_1523_ heichips25_sap3/_1524_ VPWR VGND sg13g2_and4_1
Xheichips25_sap3__3083_ heichips25_sap3/_0696_ heichips25_sap3/_1753_ heichips25_sap3/_0690_
+ heichips25_sap3/_0695_ VPWR VGND sg13g2_and3_1
Xheichips25_can_lehmann_fsm__2841__814 VPWR VGND net813 sg13g2_tiehi
XFILLER_41_795 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2034_ heichips25_sap3/net248 heichips25_sap3/_1447_ heichips25_sap3/_1440_
+ heichips25_sap3/_1455_ VPWR VGND sg13g2_a21o_1
XFILLER_13_453 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm_hold1270 heichips25_can_lehmann_fsm__2795_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1269 sg13g2_dlygate4sd3_1
XFILLER_40_272 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3985_ heichips25_sap3/net441 VGND VPWR heichips25_sap3/_0126_ heichips25_sap3__3985_/Q
+ heichips25_sap3__4009_/CLK sg13g2_dfrbpq_1
Xheichips25_sap3__2936_ heichips25_sap3/_0575_ heichips25_sap3/net276 heichips25_sap3/net211
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__2867_ heichips25_sap3/_0509_ heichips25_sap3/_0445_ heichips25_sap3/_0377_
+ heichips25_sap3/_0404_ heichips25_sap3/net154 VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2798_ heichips25_sap3/_1870_ heichips25_sap3/_0442_ heichips25_sap3/_0443_
+ VPWR VGND sg13g2_nor2_1
XFILLER_4_99 VPWR VGND sg13g2_decap_4
XFILLER_48_361 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3419_ heichips25_sap3/net121 VPWR heichips25_sap3/_1026_ VGND heichips25_sap3/net126
+ heichips25_sap3/_1025_ sg13g2_o21ai_1
XFILLER_36_567 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2640_ heichips25_can_lehmann_fsm/net468 VPWR heichips25_can_lehmann_fsm/_0786_
+ VGND heichips25_can_lehmann_fsm__2994_/Q heichips25_can_lehmann_fsm/net359 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2571_ VGND VPWR heichips25_can_lehmann_fsm/_0905_ heichips25_can_lehmann_fsm/net418
+ heichips25_can_lehmann_fsm/_0185_ heichips25_can_lehmann_fsm/_0751_ sg13g2_a21oi_1
XFILLER_32_762 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2892__712 VPWR VGND net711 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__3054_ net702 VGND VPWR heichips25_can_lehmann_fsm/_0279_
+ heichips25_can_lehmann_fsm__3054_/Q clknet_leaf_15_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2005_ heichips25_can_lehmann_fsm/net1242 heichips25_can_lehmann_fsm/net181
+ heichips25_can_lehmann_fsm/_0360_ VPWR VGND sg13g2_nor2_1
Xheichips25_can_lehmann_fsm__2907_ net681 VGND VPWR heichips25_can_lehmann_fsm/net901
+ heichips25_can_lehmann_fsm__2907_/Q clknet_leaf_12_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2838_ net530 VGND VPWR heichips25_can_lehmann_fsm/_0063_
+ heichips25_can_lehmann_fsm__2838_/Q clknet_leaf_4_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2769_ VGND VPWR heichips25_can_lehmann_fsm/_0852_ heichips25_can_lehmann_fsm/net361
+ heichips25_can_lehmann_fsm/_0284_ heichips25_can_lehmann_fsm/_0850_ sg13g2_a21oi_1
Xfanout43 uio_out_sap3\[6\] net43 VPWR VGND sg13g2_buf_2
XFILLER_23_773 VPWR VGND sg13g2_decap_4
XFILLER_10_423 VPWR VGND sg13g2_fill_2
XFILLER_6_405 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3770_ heichips25_sap3__4043_/Q heichips25_sap3__4042_/Q heichips25_sap3/_1258_
+ heichips25_sap3/_1282_ VPWR VGND sg13g2_nor3_1
Xheichips25_can_lehmann_fsm__2793__621 VPWR VGND net620 sg13g2_tiehi
Xheichips25_sap3__2721_ VGND VPWR heichips25_sap3/_0357_ heichips25_sap3/_0366_ heichips25_sap3/_0367_
+ heichips25_sap3/_0358_ sg13g2_a21oi_1
XFILLER_1_132 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2652_ VGND VPWR heichips25_sap3/net238 heichips25_sap3/_1640_ heichips25_sap3/_0319_
+ heichips25_sap3/_1784_ sg13g2_a21oi_1
Xheichips25_sap3__2583_ heichips25_sap3/_0252_ heichips25_sap3/_0253_ heichips25_sap3/_0254_
+ heichips25_sap3/_0255_ heichips25_sap3/_0256_ VPWR VGND sg13g2_and4_1
Xheichips25_can_lehmann_fsm__2869__758 VPWR VGND net757 sg13g2_tiehi
XFILLER_46_865 VPWR VGND sg13g2_decap_4
XFILLER_45_331 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3204_ heichips25_sap3/_0817_ heichips25_sap3__3966_/Q heichips25_sap3/net144
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__3135_ VPWR heichips25_sap3/_0748_ heichips25_sap3/_0747_ VGND sg13g2_inv_1
XFILLER_33_548 VPWR VGND sg13g2_decap_8
XFILLER_33_559 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3066_ heichips25_sap3/_0679_ heichips25_sap3/_0676_ heichips25_sap3/_0677_
+ VPWR VGND sg13g2_nand2_1
XFILLER_20_209 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2017_ VGND VPWR heichips25_sap3/_1438_ heichips25_sap3/net261 heichips25_sap3/net262
+ sg13g2_or2_1
XFILLER_9_243 VPWR VGND sg13g2_fill_2
XFILLER_9_254 VPWR VGND sg13g2_decap_8
Xclkload13 clkload13/Y clknet_leaf_8_clk VPWR VGND sg13g2_inv_2
Xclkload24 VPWR clkload24/Y clkload24/A VGND sg13g2_inv_1
Xheichips25_sap3__3968_ heichips25_sap3/net441 VGND VPWR heichips25_sap3/_0109_ heichips25_sap3__3968_/Q
+ heichips25_sap3__4016_/CLK sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm_fanout308 heichips25_can_lehmann_fsm/net309 heichips25_can_lehmann_fsm/net308
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout319 heichips25_can_lehmann_fsm/net320 heichips25_can_lehmann_fsm/net319
+ VPWR VGND sg13g2_buf_1
Xheichips25_sap3__2919_ heichips25_sap3/net69 heichips25_sap3/_0538_ heichips25_sap3/_0558_
+ heichips25_sap3/_0559_ VPWR VGND sg13g2_nor3_1
Xheichips25_sap3__3899_ heichips25_sap3/net447 VGND VPWR heichips25_sap3/_0040_ heichips25_sap3__3899_/Q
+ heichips25_sap3__4003_/CLK sg13g2_dfrbpq_1
XFILLER_49_670 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2623_ VGND VPWR heichips25_can_lehmann_fsm/_0892_ heichips25_can_lehmann_fsm/net416
+ heichips25_can_lehmann_fsm/_0211_ heichips25_can_lehmann_fsm/_0777_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2554_ heichips25_can_lehmann_fsm/net494 VPWR heichips25_can_lehmann_fsm/_0743_
+ VGND heichips25_can_lehmann_fsm/net1082 heichips25_can_lehmann_fsm/net407 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2485_ VGND VPWR heichips25_can_lehmann_fsm/_0926_ heichips25_can_lehmann_fsm/net368
+ heichips25_can_lehmann_fsm/_0142_ heichips25_can_lehmann_fsm/_0708_ sg13g2_a21oi_1
Xclkload7 VPWR clkload7/Y clknet_leaf_5_clk VGND sg13g2_inv_1
XFILLER_3_419 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__3037_ net806 VGND VPWR heichips25_can_lehmann_fsm/_0262_
+ heichips25_can_lehmann_fsm__3037_/Q clknet_leaf_20_clk sg13g2_dfrbpq_1
XFILLER_8_1024 VPWR VGND sg13g2_decap_4
XFILLER_46_117 VPWR VGND sg13g2_fill_2
XFILLER_42_367 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_hold942 heichips25_can_lehmann_fsm__2856_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net941 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold920 heichips25_can_lehmann_fsm/_0216_ VPWR VGND heichips25_can_lehmann_fsm/net919
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold953 heichips25_can_lehmann_fsm/_0256_ VPWR VGND heichips25_can_lehmann_fsm/net952
+ sg13g2_dlygate4sd3_1
XFILLER_24_63 VPWR VGND sg13g2_decap_8
XFILLER_24_74 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm_hold931 heichips25_can_lehmann_fsm__2976_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net930 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold975 heichips25_can_lehmann_fsm__2842_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net974 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold964 heichips25_can_lehmann_fsm__2988_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net963 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__2940__576 VPWR VGND net575 sg13g2_tiehi
Xheichips25_can_lehmann_fsm_hold986 heichips25_can_lehmann_fsm__2983_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net985 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold997 heichips25_can_lehmann_fsm__2903_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net996 sg13g2_dlygate4sd3_1
Xheichips25_sap3__3822_ heichips25_sap3/_1328_ heichips25_sap3/net292 heichips25_sap3__3961_/Q
+ heichips25_sap3/_1259_ heichips25_sap3__3985_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3753_ heichips25_sap3__4040_/Q heichips25_sap3__4041_/Q heichips25_sap3/_1264_
+ heichips25_sap3/_1265_ VPWR VGND sg13g2_nor3_1
Xheichips25_sap3__2704_ heichips25_sap3__3921_/Q heichips25_sap3/net276 heichips25_sap3/_0350_
+ VPWR VGND sg13g2_xor2_1
Xheichips25_sap3__3684_ VPWR heichips25_sap3/_0144_ heichips25_sap3/_1224_ VGND sg13g2_inv_1
XFILLER_49_82 VPWR VGND sg13g2_decap_8
XFILLER_49_60 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2635_ VGND VPWR heichips25_sap3/_0297_ heichips25_sap3/_0301_ heichips25_sap3/_0302_
+ heichips25_sap3/net244 sg13g2_a21oi_1
X_21_ net522 net47 net505 net34 VPWR VGND sg13g2_mux2_1
Xheichips25_sap3__2566_ VGND VPWR heichips25_sap3/_0237_ heichips25_sap3/_0240_ heichips25_sap3/_0241_
+ heichips25_sap3/net66 sg13g2_a21oi_1
Xheichips25_sap3__2497_ heichips25_sap3/_1910_ heichips25_sap3__3893_/Q heichips25_sap3/_1788_
+ VPWR VGND sg13g2_nand2_1
XFILLER_18_364 VPWR VGND sg13g2_fill_1
XFILLER_18_375 VPWR VGND sg13g2_fill_2
XFILLER_33_334 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3118_ VPWR VGND heichips25_sap3/_1363_ heichips25_sap3/_0730_ heichips25_sap3/_0654_
+ heichips25_sap3/net247 heichips25_sap3/_0731_ heichips25_sap3/net246 sg13g2_a221oi_1
Xheichips25_sap3__3049_ heichips25_sap3/_1455_ heichips25_sap3/_1465_ heichips25_sap3/_0661_
+ heichips25_sap3/_0662_ VPWR VGND sg13g2_nor3_1
Xheichips25_can_lehmann_fsm__2270_ VGND VPWR heichips25_can_lehmann_fsm/net207 heichips25_can_lehmann_fsm/_0585_
+ heichips25_can_lehmann_fsm/_0049_ heichips25_can_lehmann_fsm/_0586_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__1985_ VPWR VGND heichips25_can_lehmann_fsm/net1234 heichips25_can_lehmann_fsm/net194
+ heichips25_can_lehmann_fsm/net189 heichips25_can_lehmann_fsm__2782_/Q heichips25_can_lehmann_fsm/_0343_
+ heichips25_can_lehmann_fsm/net197 sg13g2_a221oi_1
XFILLER_25_813 VPWR VGND sg13g2_decap_8
XFILLER_24_356 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2606_ heichips25_can_lehmann_fsm/net491 VPWR heichips25_can_lehmann_fsm/_0769_
+ VGND heichips25_can_lehmann_fsm/net897 heichips25_can_lehmann_fsm/net422 sg13g2_o21ai_1
XFILLER_25_879 VPWR VGND sg13g2_fill_2
XFILLER_40_849 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2537_ VGND VPWR heichips25_can_lehmann_fsm/_0913_ heichips25_can_lehmann_fsm/net357
+ heichips25_can_lehmann_fsm/_0168_ heichips25_can_lehmann_fsm/_0734_ sg13g2_a21oi_1
XFILLER_20_551 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2468_ heichips25_can_lehmann_fsm/net498 VPWR heichips25_can_lehmann_fsm/_0700_
+ VGND heichips25_can_lehmann_fsm/net903 heichips25_can_lehmann_fsm/net384 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2399_ VGND VPWR heichips25_can_lehmann_fsm/_0951_ heichips25_can_lehmann_fsm/net355
+ heichips25_can_lehmann_fsm/_0099_ heichips25_can_lehmann_fsm/_0665_ sg13g2_a21oi_1
XFILLER_3_216 VPWR VGND sg13g2_fill_2
XFILLER_10_10 VPWR VGND sg13g2_fill_1
XFILLER_10_43 VPWR VGND sg13g2_decap_8
XFILLER_0_901 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2420_ heichips25_sap3/_1837_ heichips25_sap3/net78 heichips25_sap3__4024_/Q
+ heichips25_sap3/net86 heichips25_sap3__3960_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_0_978 VPWR VGND sg13g2_decap_8
XFILLER_19_52 VPWR VGND sg13g2_decap_8
XFILLER_19_74 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2351_ heichips25_sap3/_1454_ heichips25_sap3/net226 heichips25_sap3/_1613_
+ heichips25_sap3/_1772_ VPWR VGND sg13g2_nor3_1
Xheichips25_sap3__2282_ heichips25_sap3/_1703_ heichips25_sap3/_1629_ heichips25_sap3/_1702_
+ VPWR VGND sg13g2_nand2_1
XFILLER_16_835 VPWR VGND sg13g2_decap_8
XFILLER_43_654 VPWR VGND sg13g2_decap_8
XFILLER_42_120 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__4021_ heichips25_sap3/net449 VGND VPWR heichips25_sap3/_0162_ heichips25_sap3__4021_/Q
+ heichips25_sap3__4021_/CLK sg13g2_dfrbpq_1
XFILLER_35_73 VPWR VGND sg13g2_fill_2
XFILLER_31_805 VPWR VGND sg13g2_fill_2
XFILLER_31_816 VPWR VGND sg13g2_fill_1
XFILLER_43_698 VPWR VGND sg13g2_fill_2
XFILLER_31_838 VPWR VGND sg13g2_fill_1
XFILLER_30_348 VPWR VGND sg13g2_decap_8
XFILLER_7_511 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__1997_ VPWR heichips25_sap3/_1423_ heichips25_sap3__3986_/Q VGND
+ sg13g2_inv_1
Xheichips25_sap3__3805_ heichips25_sap3/_1313_ heichips25_sap3/_1281_ heichips25_sap3__4015_/Q
+ heichips25_sap3/_1259_ heichips25_sap3__3983_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3736_ VPWR VGND heichips25_sap3/_1252_ heichips25_sap3/_1251_ heichips25_sap3/_0290_
+ heichips25_sap3/_1360_ heichips25_sap3/_1253_ heichips25_sap3__4032_/Q sg13g2_a221oi_1
Xheichips25_sap3__3667_ heichips25_sap3/net111 heichips25_sap3__3999_/Q heichips25_sap3/_1211_
+ heichips25_sap3/_0140_ VPWR VGND sg13g2_a21o_1
XFILLER_3_783 VPWR VGND sg13g2_decap_8
XFILLER_2_260 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2618_ heichips25_sap3/_0286_ heichips25_sap3/_0287_ heichips25_sap3/_0288_
+ VPWR VGND sg13g2_nor2b_1
Xheichips25_sap3__3598_ VGND VPWR heichips25_sap3/net137 heichips25_sap3/net131 heichips25_sap3/_1171_
+ heichips25_sap3/net139 sg13g2_a21oi_1
X_04_ net507 net2 _00_ VPWR VGND sg13g2_nor2b_1
Xheichips25_sap3__2549_ heichips25_sap3/_0033_ heichips25_sap3/_1925_ heichips25_sap3/_0224_
+ VPWR VGND sg13g2_nand2_1
XFILLER_47_971 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1770_ heichips25_can_lehmann_fsm/_1086_ heichips25_can_lehmann_fsm/net310
+ heichips25_can_lehmann_fsm__3014_/Q heichips25_can_lehmann_fsm/net313 heichips25_can_lehmann_fsm__2918_/Q
+ VPWR VGND sg13g2_a22oi_1
XFILLER_18_150 VPWR VGND sg13g2_decap_8
XFILLER_18_161 VPWR VGND sg13g2_decap_8
XFILLER_33_153 VPWR VGND sg13g2_decap_8
XFILLER_21_304 VPWR VGND sg13g2_decap_8
XFILLER_21_326 VPWR VGND sg13g2_fill_2
XFILLER_21_348 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2322_ heichips25_can_lehmann_fsm/net471 VPWR heichips25_can_lehmann_fsm/_0627_
+ VGND heichips25_can_lehmann_fsm/net1136 heichips25_can_lehmann_fsm/net403 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2253_ heichips25_can_lehmann_fsm/net327 VPWR heichips25_can_lehmann_fsm/_0573_
+ VGND heichips25_can_lehmann_fsm/net1173 heichips25_can_lehmann_fsm/net206 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2184_ VGND VPWR heichips25_can_lehmann_fsm/_0516_ heichips25_can_lehmann_fsm/_0517_
+ heichips25_can_lehmann_fsm/_0031_ heichips25_can_lehmann_fsm/_0518_ sg13g2_a21oi_1
XFILLER_29_415 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1968_ heichips25_can_lehmann_fsm__2782_/Q heichips25_can_lehmann_fsm/_0304_
+ heichips25_can_lehmann_fsm/_0328_ VPWR VGND sg13g2_and2_1
XFILLER_16_109 VPWR VGND sg13g2_fill_1
XFILLER_25_621 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1899_ VGND VPWR heichips25_can_lehmann_fsm__2905_/Q heichips25_can_lehmann_fsm/net297
+ heichips25_can_lehmann_fsm/_1212_ heichips25_can_lehmann_fsm/_1211_ sg13g2_a21oi_1
Xheichips25_sap3_hold1121 heichips25_sap3__4034_/Q VPWR VGND heichips25_sap3/net1120
+ sg13g2_dlygate4sd3_1
Xheichips25_sap3_hold1132 heichips25_sap3/_0291_ VPWR VGND heichips25_sap3/net1131
+ sg13g2_dlygate4sd3_1
XFILLER_25_698 VPWR VGND sg13g2_fill_2
Xheichips25_sap3_hold1198 heichips25_sap3__4040_/Q VPWR VGND heichips25_sap3/net1197
+ sg13g2_dlygate4sd3_1
XFILLER_40_668 VPWR VGND sg13g2_fill_1
XFILLER_20_381 VPWR VGND sg13g2_fill_2
XFILLER_4_525 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_fanout491 heichips25_can_lehmann_fsm/net496 heichips25_can_lehmann_fsm/net491
+ VPWR VGND sg13g2_buf_1
Xheichips25_sap3__3521_ heichips25_sap3/_1114_ heichips25_sap3/_0749_ heichips25_sap3/_0977_
+ VPWR VGND sg13g2_nand2b_1
Xheichips25_can_lehmann_fsm_fanout480 heichips25_can_lehmann_fsm/net481 heichips25_can_lehmann_fsm/net480
+ VPWR VGND sg13g2_buf_1
Xheichips25_sap3__3452_ heichips25_sap3/_1057_ heichips25_sap3/net60 heichips25_sap3/net99
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__3383_ heichips25_sap3/_0991_ heichips25_sap3/_0985_ heichips25_sap3/_0990_
+ heichips25_sap3/net124 heichips25_sap3/_1404_ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2403_ VPWR VGND heichips25_sap3__3961_/Q heichips25_sap3/_1821_
+ heichips25_sap3/net85 heichips25_sap3__3953_/Q heichips25_sap3/_1822_ heichips25_sap3/net87
+ sg13g2_a221oi_1
XFILLER_47_289 VPWR VGND sg13g2_fill_1
XFILLER_35_418 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2334_ heichips25_sap3/net242 heichips25_sap3/_1549_ heichips25_sap3/net266
+ heichips25_sap3/_1755_ VPWR VGND sg13g2_nand3_1
XFILLER_29_960 VPWR VGND sg13g2_fill_2
XFILLER_46_72 VPWR VGND sg13g2_decap_8
XFILLER_28_470 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2265_ VGND VPWR heichips25_sap3/net236 heichips25_sap3/_1474_ heichips25_sap3/_1686_
+ heichips25_sap3/net245 sg13g2_a21oi_1
Xheichips25_sap3__4004_ heichips25_sap3/net436 VGND VPWR heichips25_sap3/_0145_ heichips25_sap3__4004_/Q
+ heichips25_sap3__4005_/CLK sg13g2_dfrbpq_1
Xheichips25_sap3__2196_ heichips25_sap3/_1615_ heichips25_sap3/_1616_ heichips25_sap3/_1617_
+ VPWR VGND sg13g2_nor2_1
XFILLER_15_164 VPWR VGND sg13g2_decap_8
XFILLER_7_44 VPWR VGND sg13g2_fill_1
XFILLER_11_392 VPWR VGND sg13g2_fill_1
XFILLER_7_363 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3719_ heichips25_sap3__4020_/Q heichips25_sap3/_1175_ heichips25_sap3/net117
+ heichips25_sap3/_0161_ VPWR VGND sg13g2_mux2_1
Xheichips25_can_lehmann_fsm__2940_ net575 VGND VPWR heichips25_can_lehmann_fsm/_0165_
+ heichips25_can_lehmann_fsm__2940_/Q clknet_leaf_18_clk sg13g2_dfrbpq_1
XFILLER_39_779 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2871_ net753 VGND VPWR heichips25_can_lehmann_fsm/_0096_
+ heichips25_can_lehmann_fsm__2871_/Q clknet_leaf_20_clk sg13g2_dfrbpq_1
XFILLER_26_429 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1822_ VGND VPWR heichips25_can_lehmann_fsm/_1136_ heichips25_can_lehmann_fsm/_1137_
+ heichips25_can_lehmann_fsm/_1138_ heichips25_can_lehmann_fsm/_1133_ sg13g2_a21oi_1
XFILLER_35_941 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1753_ heichips25_can_lehmann_fsm__2790_/Q heichips25_can_lehmann_fsm/_1072_
+ heichips25_can_lehmann_fsm/_1073_ VPWR VGND sg13g2_nor2_1
Xheichips25_can_lehmann_fsm__1684_ VGND VPWR heichips25_can_lehmann_fsm__2945_/Q heichips25_can_lehmann_fsm/net305
+ heichips25_can_lehmann_fsm/_1008_ heichips25_can_lehmann_fsm/net300 sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__3025__683 VPWR VGND net682 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2305_ heichips25_can_lehmann_fsm/net327 VPWR heichips25_can_lehmann_fsm/_0615_
+ VGND heichips25_can_lehmann_fsm/net1158 heichips25_can_lehmann_fsm/net209 sg13g2_o21ai_1
Xclkbuf_5_28__f_heichips25_sap3\_sap_3_inst.alu_inst.clk heichips25_sap3__3990_/CLK
+ clknet_4_14_0_heichips25_sap3\/sap_3_inst.alu_inst.clk VPWR VGND sg13g2_buf_16
Xheichips25_can_lehmann_fsm__2236_ VGND VPWR heichips25_can_lehmann_fsm/net857 heichips25_can_lehmann_fsm/net170
+ heichips25_can_lehmann_fsm/_0559_ heichips25_can_lehmann_fsm/_0558_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2167_ heichips25_can_lehmann_fsm/net325 VPWR heichips25_can_lehmann_fsm/_0505_
+ VGND heichips25_can_lehmann_fsm/net1233 heichips25_can_lehmann_fsm/net160 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2098_ heichips25_can_lehmann_fsm/_0439_ heichips25_can_lehmann_fsm/net196
+ net17 heichips25_can_lehmann_fsm/net199 heichips25_can_lehmann_fsm/net1270 VPWR
+ VGND sg13g2_a22oi_1
XFILLER_18_908 VPWR VGND sg13g2_fill_2
XFILLER_18_919 VPWR VGND sg13g2_fill_1
XFILLER_29_278 VPWR VGND sg13g2_fill_1
XFILLER_17_429 VPWR VGND sg13g2_fill_1
XFILLER_26_941 VPWR VGND sg13g2_fill_1
Xheichips25_sap3_fanout340 heichips25_sap3/_0008_ heichips25_sap3/net340 VPWR VGND
+ sg13g2_buf_1
XFILLER_41_933 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2050_ heichips25_sap3/_1471_ heichips25_sap3/_1469_ heichips25_sap3/_1470_
+ VPWR VGND sg13g2_nand2b_1
XFILLER_25_484 VPWR VGND sg13g2_fill_1
XFILLER_9_617 VPWR VGND sg13g2_decap_4
XFILLER_9_639 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2952_ heichips25_sap3/_0590_ heichips25_sap3/_0449_ heichips25_sap3/_0348_
+ VPWR VGND sg13g2_nand2b_1
Xheichips25_sap3__2883_ heichips25_sap3/_0406_ heichips25_sap3/_0405_ heichips25_sap3/_0524_
+ VPWR VGND sg13g2_xor2_1
XFILLER_10_1021 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3504_ heichips25_sap3/_0089_ heichips25_sap3/_1095_ heichips25_sap3/_1099_
+ heichips25_sap3/net106 heichips25_sap3/_1391_ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3435_ heichips25_sap3/_1040_ VPWR heichips25_sap3/_1041_ VGND heichips25_sap3/_0720_
+ heichips25_sap3/_1037_ sg13g2_o21ai_1
Xclkbuf_4_2_0_heichips25_sap3\_sap_3_inst.alu_inst.clk clknet_0_heichips25_sap3\/sap_3_inst.alu_inst.clk
+ clknet_4_2_0_heichips25_sap3\/sap_3_inst.alu_inst.clk VPWR VGND sg13g2_buf_8
Xheichips25_sap3__3366_ heichips25_sap3/_0971_ heichips25_sap3/net124 heichips25_sap3/_0974_
+ heichips25_sap3/_0975_ VPWR VGND sg13g2_a21o_1
XFILLER_17_941 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2317_ heichips25_sap3/_1738_ heichips25_sap3/net85 heichips25_sap3__3954_/Q
+ heichips25_sap3/net87 heichips25_sap3__3946_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3297_ heichips25_sap3/net48 heichips25_sap3/net51 heichips25_sap3/net59
+ heichips25_sap3/_0909_ VPWR VGND sg13g2_nand3_1
XFILLER_44_782 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2248_ heichips25_sap3/net223 heichips25_sap3/_1668_ heichips25_sap3/net240
+ heichips25_sap3/_1669_ VPWR VGND sg13g2_nand3_1
XFILLER_16_462 VPWR VGND sg13g2_fill_1
XFILLER_31_410 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2179_ heichips25_sap3/_1523_ heichips25_sap3/_1561_ heichips25_sap3/_1600_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_can_lehmann_fsm__2879__738 VPWR VGND net737 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2994__642 VPWR VGND net641 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2021_ heichips25_can_lehmann_fsm/net1246 VPWR heichips25_can_lehmann_fsm/_0373_
+ VGND heichips25_can_lehmann_fsm__2788_/Q heichips25_can_lehmann_fsm/_1070_ sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2923_ net643 VGND VPWR heichips25_can_lehmann_fsm/_0148_
+ heichips25_can_lehmann_fsm__2923_/Q clknet_leaf_0_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2854_ net787 VGND VPWR heichips25_can_lehmann_fsm/net899
+ heichips25_can_lehmann_fsm__2854_/Q clknet_leaf_9_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2785_ net636 VGND VPWR heichips25_can_lehmann_fsm/net1252
+ heichips25_can_lehmann_fsm__2785_/Q clknet_leaf_5_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1805_ heichips25_can_lehmann_fsm/_1117_ heichips25_can_lehmann_fsm/_1118_
+ heichips25_can_lehmann_fsm/_1119_ heichips25_can_lehmann_fsm/_1120_ heichips25_can_lehmann_fsm/_1121_
+ VPWR VGND sg13g2_and4_1
Xheichips25_can_lehmann_fsm__1736_ heichips25_can_lehmann_fsm__2797_/Q heichips25_can_lehmann_fsm/net346
+ heichips25_can_lehmann_fsm/net347 heichips25_can_lehmann_fsm__2794_/Q heichips25_can_lehmann_fsm/_1056_
+ VPWR VGND sg13g2_or4_1
Xheichips25_can_lehmann_fsm__1667_ heichips25_can_lehmann_fsm/net353 heichips25_can_lehmann_fsm/net350
+ heichips25_can_lehmann_fsm/_0991_ VPWR VGND heichips25_can_lehmann_fsm/net351 sg13g2_nand3b_1
Xheichips25_can_lehmann_fsm__1598_ VPWR heichips25_can_lehmann_fsm/_0922_ heichips25_can_lehmann_fsm/net1047
+ VGND sg13g2_inv_1
XFILLER_5_119 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2219_ heichips25_can_lehmann_fsm/net329 VPWR heichips25_can_lehmann_fsm/_0546_
+ VGND heichips25_can_lehmann_fsm/net1231 heichips25_can_lehmann_fsm/net162 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2936__592 VPWR VGND net591 sg13g2_tiehi
Xheichips25_sap3__3220_ heichips25_sap3/_0833_ heichips25_sap3/net138 heichips25_sap3__3981_/Q
+ heichips25_sap3/net140 heichips25_sap3__3989_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_45_524 VPWR VGND sg13g2_fill_2
XFILLER_45_513 VPWR VGND sg13g2_decap_4
XFILLER_27_30 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3151_ VPWR heichips25_sap3/_0764_ heichips25_sap3/net104 VGND sg13g2_inv_1
XFILLER_27_96 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2102_ heichips25_sap3/net242 heichips25_sap3/_1522_ heichips25_sap3/_1523_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__3082_ heichips25_sap3/_0694_ VPWR heichips25_sap3/_0695_ VGND heichips25_sap3/net220
+ heichips25_sap3/_0693_ sg13g2_o21ai_1
XFILLER_32_218 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2033_ heichips25_sap3/_1454_ heichips25_sap3/_1443_ heichips25_sap3/_1449_
+ VPWR VGND sg13g2_nand2_1
XFILLER_25_281 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm_hold1260 heichips25_can_lehmann_fsm__2788_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1259 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1271 heichips25_can_lehmann_fsm__2799_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1270 sg13g2_dlygate4sd3_1
XFILLER_9_447 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3984_ heichips25_sap3/net441 VGND VPWR heichips25_sap3/_0125_ heichips25_sap3__3984_/Q
+ clkload20/A sg13g2_dfrbpq_1
Xheichips25_sap3__2935_ heichips25_sap3/net65 heichips25_sap3/_0565_ heichips25_sap3/_0573_
+ heichips25_sap3/_0574_ VPWR VGND sg13g2_nor3_1
XFILLER_4_130 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2866_ heichips25_sap3/_0508_ heichips25_sap3/_0500_ heichips25_sap3/_0338_
+ heichips25_sap3/_0498_ heichips25_sap3/_0340_ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2797_ heichips25_sap3/_1880_ heichips25_sap3/_1881_ heichips25_sap3/_1884_
+ heichips25_sap3/net168 heichips25_sap3/_0442_ VPWR VGND sg13g2_and4_1
XFILLER_4_67 VPWR VGND sg13g2_fill_1
X_21__523 VPWR VGND net522 sg13g2_tielo
XFILLER_49_874 VPWR VGND sg13g2_fill_1
XFILLER_48_373 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3418_ heichips25_sap3/_1025_ heichips25_sap3/_0794_ heichips25_sap3/_0856_
+ VPWR VGND sg13g2_xnor2_1
XFILLER_36_579 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3349_ heichips25_sap3/_0075_ heichips25_sap3/_0950_ heichips25_sap3/_0958_
+ heichips25_sap3/net55 heichips25_sap3/_1368_ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2570_ heichips25_can_lehmann_fsm/net487 VPWR heichips25_can_lehmann_fsm/_0751_
+ VGND heichips25_can_lehmann_fsm__2960_/Q heichips25_can_lehmann_fsm/net418 sg13g2_o21ai_1
XFILLER_31_295 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__3053_ net734 VGND VPWR heichips25_can_lehmann_fsm/net1052
+ heichips25_can_lehmann_fsm__3053_/Q clknet_leaf_12_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2004_ heichips25_can_lehmann_fsm/_0359_ heichips25_can_lehmann_fsm/net184
+ heichips25_can_lehmann_fsm/_0358_ heichips25_can_lehmann_fsm/net197 heichips25_can_lehmann_fsm__2785_/Q
+ VPWR VGND sg13g2_a22oi_1
XFILLER_39_373 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2906_ net683 VGND VPWR heichips25_can_lehmann_fsm/_0131_
+ heichips25_can_lehmann_fsm__2906_/Q clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_27_524 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2837_ net532 VGND VPWR heichips25_can_lehmann_fsm/net896
+ heichips25_can_lehmann_fsm__2837_/Q clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_14_218 VPWR VGND sg13g2_decap_8
XFILLER_27_579 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2768_ heichips25_can_lehmann_fsm/net480 VPWR heichips25_can_lehmann_fsm/_0850_
+ VGND heichips25_can_lehmann_fsm__3058_/Q heichips25_can_lehmann_fsm/net361 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2699_ VGND VPWR heichips25_can_lehmann_fsm/_0870_ heichips25_can_lehmann_fsm/net382
+ heichips25_can_lehmann_fsm/_0249_ heichips25_can_lehmann_fsm/_0815_ sg13g2_a21oi_1
Xfanout44 uio_out_sap3\[2\] net44 VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm__1719_ heichips25_can_lehmann_fsm/_1041_ heichips25_can_lehmann_fsm/_1034_
+ heichips25_can_lehmann_fsm/net1213 heichips25_can_lehmann_fsm/_1029_ heichips25_can_lehmann_fsm/_1016_
+ VPWR VGND sg13g2_a22oi_1
XFILLER_13_21 VPWR VGND sg13g2_decap_8
XFILLER_10_446 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2720_ VGND VPWR heichips25_sap3/_0361_ heichips25_sap3/_0365_ heichips25_sap3/_0366_
+ heichips25_sap3/_0360_ sg13g2_a21oi_1
Xheichips25_sap3__2651_ heichips25_sap3/_1641_ VPWR heichips25_sap3/_0318_ VGND heichips25_sap3/_0311_
+ heichips25_sap3/_0317_ sg13g2_o21ai_1
XFILLER_49_137 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2582_ heichips25_sap3/_0255_ heichips25_sap3/net76 heichips25_sap3__3981_/Q
+ heichips25_sap3/net78 heichips25_sap3__4013_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_45_354 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3203_ heichips25_sap3/_0816_ heichips25_sap3/net105 heichips25_sap3__3950_/Q
+ heichips25_sap3/net108 heichips25_sap3__3958_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_18_579 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3134_ VGND VPWR heichips25_sap3/_0737_ heichips25_sap3/_0746_ heichips25_sap3/_0747_
+ heichips25_sap3/net123 sg13g2_a21oi_1
Xheichips25_sap3__3065_ heichips25_sap3/_0676_ heichips25_sap3/_0677_ heichips25_sap3/_0678_
+ VPWR VGND sg13g2_and2_1
Xheichips25_sap3__2016_ VGND VPWR heichips25_sap3/_1437_ heichips25_sap3/net264 heichips25_sap3/net267
+ sg13g2_or2_1
XFILLER_13_273 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_hold1090 heichips25_can_lehmann_fsm/_0066_ VPWR VGND heichips25_can_lehmann_fsm/net1089
+ sg13g2_dlygate4sd3_1
XFILLER_13_295 VPWR VGND sg13g2_fill_1
Xclkload14 clknet_leaf_9_clk clkload14/X VPWR VGND sg13g2_buf_8
Xclkload25 VPWR clkload25/Y clkload25/A VGND sg13g2_inv_1
Xheichips25_sap3__3967_ heichips25_sap3/net443 VGND VPWR heichips25_sap3/_0108_ heichips25_sap3__3967_/Q
+ heichips25_sap3__4009_/CLK sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm_fanout309 heichips25_can_lehmann_fsm/_0997_ heichips25_can_lehmann_fsm/net309
+ VPWR VGND sg13g2_buf_1
Xheichips25_sap3__2918_ VPWR VGND heichips25_sap3/_0557_ heichips25_sap3/net157 heichips25_sap3/_0556_
+ heichips25_sap3__3912_/Q heichips25_sap3/_0558_ heichips25_sap3/net203 sg13g2_a221oi_1
Xheichips25_sap3__3898_ heichips25_sap3/net450 VGND VPWR heichips25_sap3/_0039_ heichips25_sap3__3898_/Q
+ clkload23/A sg13g2_dfrbpq_1
Xheichips25_sap3__2849_ heichips25_sap3/_0481_ heichips25_sap3/_0488_ heichips25_sap3/_0480_
+ heichips25_sap3/_0492_ VPWR VGND heichips25_sap3/_0491_ sg13g2_nand4_1
XFILLER_36_332 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2622_ heichips25_can_lehmann_fsm/net484 VPWR heichips25_can_lehmann_fsm/_0777_
+ VGND heichips25_can_lehmann_fsm__2986_/Q heichips25_can_lehmann_fsm/net416 sg13g2_o21ai_1
XFILLER_24_538 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2553_ VGND VPWR heichips25_can_lehmann_fsm/_0909_ heichips25_can_lehmann_fsm/net367
+ heichips25_can_lehmann_fsm/_0176_ heichips25_can_lehmann_fsm/_0742_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2484_ heichips25_can_lehmann_fsm/net477 VPWR heichips25_can_lehmann_fsm/_0708_
+ VGND heichips25_can_lehmann_fsm/net1135 heichips25_can_lehmann_fsm/net368 sg13g2_o21ai_1
Xclkload8 clkload8/Y clknet_leaf_7_clk VPWR VGND sg13g2_inv_2
Xheichips25_can_lehmann_fsm__3036_ net533 VGND VPWR heichips25_can_lehmann_fsm/_0261_
+ heichips25_can_lehmann_fsm__3036_/Q clknet_leaf_20_clk sg13g2_dfrbpq_1
XFILLER_28_800 VPWR VGND sg13g2_fill_2
XFILLER_39_170 VPWR VGND sg13g2_decap_4
XFILLER_27_332 VPWR VGND sg13g2_decap_8
XFILLER_28_877 VPWR VGND sg13g2_decap_4
XFILLER_15_527 VPWR VGND sg13g2_fill_2
XFILLER_27_354 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm_hold910 heichips25_can_lehmann_fsm__2909_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net909 sg13g2_dlygate4sd3_1
XFILLER_30_519 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm_hold943 heichips25_can_lehmann_fsm__2859_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net942 sg13g2_dlygate4sd3_1
XFILLER_11_711 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm_hold932 heichips25_can_lehmann_fsm__3005_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net931 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold921 heichips25_can_lehmann_fsm__3004_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net920 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__2905__686 VPWR VGND net685 sg13g2_tiehi
XFILLER_7_715 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm_hold965 heichips25_can_lehmann_fsm__2992_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net964 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold976 heichips25_can_lehmann_fsm__2912_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net975 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold998 heichips25_can_lehmann_fsm/_0129_ VPWR VGND heichips25_can_lehmann_fsm/net997
+ sg13g2_dlygate4sd3_1
XFILLER_6_225 VPWR VGND sg13g2_decap_8
XFILLER_6_214 VPWR VGND sg13g2_fill_2
XFILLER_10_276 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm_hold987 heichips25_can_lehmann_fsm/_0208_ VPWR VGND heichips25_can_lehmann_fsm/net986
+ sg13g2_dlygate4sd3_1
Xheichips25_sap3__3821_ VGND VPWR heichips25_sap3__4025_/Q heichips25_sap3/_1270_
+ heichips25_sap3/_1327_ heichips25_sap3/net291 sg13g2_a21oi_1
XFILLER_6_247 VPWR VGND sg13g2_decap_4
XFILLER_10_287 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3752_ heichips25_sap3/_1264_ heichips25_sap3__4043_/Q heichips25_sap3__4042_/Q
+ VPWR VGND sg13g2_nand2b_1
Xheichips25_sap3__2703_ heichips25_sap3/_1384_ heichips25_sap3/_1398_ heichips25_sap3/_0349_
+ VPWR VGND sg13g2_nor2_1
XFILLER_3_998 VPWR VGND sg13g2_decap_8
XFILLER_2_475 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3683_ heichips25_sap3/_1224_ heichips25_sap3/_1056_ heichips25_sap3/_1223_
+ heichips25_sap3/net113 heichips25_sap3__4003_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2634_ heichips25_sap3/_1568_ VPWR heichips25_sap3/_0301_ VGND heichips25_sap3/_1491_
+ heichips25_sap3/_1494_ sg13g2_o21ai_1
X_20_ net521 net43 net504 net33 VPWR VGND sg13g2_mux2_1
Xheichips25_sap3__2565_ heichips25_sap3/_0235_ heichips25_sap3/_0236_ heichips25_sap3/_0238_
+ heichips25_sap3/_0239_ heichips25_sap3/_0240_ VPWR VGND sg13g2_and4_1
XFILLER_1_68 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2496_ heichips25_sap3/_1909_ net4 heichips25_sap3/_1770_ VPWR VGND
+ sg13g2_nand2_1
XFILLER_46_663 VPWR VGND sg13g2_fill_1
XFILLER_34_825 VPWR VGND sg13g2_decap_8
XFILLER_45_184 VPWR VGND sg13g2_fill_2
XFILLER_18_387 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3117_ VGND VPWR heichips25_sap3/_0721_ heichips25_sap3/_0729_ heichips25_sap3/_0730_
+ heichips25_sap3/_0313_ sg13g2_a21oi_1
Xheichips25_sap3__3048_ VGND VPWR heichips25_sap3/net227 heichips25_sap3/_1644_ heichips25_sap3/_0661_
+ heichips25_sap3/net241 sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2806__595 VPWR VGND net594 sg13g2_tiehi
XFILLER_39_0 VPWR VGND sg13g2_fill_1
Xinput1 ena net1 VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm__1984_ heichips25_can_lehmann_fsm/net344 heichips25_can_lehmann_fsm/net193
+ heichips25_can_lehmann_fsm/_0342_ VPWR VGND sg13g2_nor2b_1
XFILLER_24_324 VPWR VGND sg13g2_fill_2
XFILLER_40_817 VPWR VGND sg13g2_fill_1
XFILLER_24_346 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2605_ VGND VPWR heichips25_can_lehmann_fsm/_0896_ heichips25_can_lehmann_fsm/net380
+ heichips25_can_lehmann_fsm/_0202_ heichips25_can_lehmann_fsm/_0768_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2536_ heichips25_can_lehmann_fsm/net476 VPWR heichips25_can_lehmann_fsm/_0734_
+ VGND heichips25_can_lehmann_fsm__2942_/Q heichips25_can_lehmann_fsm/net358 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2467_ VGND VPWR heichips25_can_lehmann_fsm/_0931_ heichips25_can_lehmann_fsm/net426
+ heichips25_can_lehmann_fsm/_0133_ heichips25_can_lehmann_fsm/_0699_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2398_ heichips25_can_lehmann_fsm/net470 VPWR heichips25_can_lehmann_fsm/_0665_
+ VGND heichips25_can_lehmann_fsm/net1080 heichips25_can_lehmann_fsm/net355 sg13g2_o21ai_1
XFILLER_10_88 VPWR VGND sg13g2_decap_8
XFILLER_0_957 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__3019_ net730 VGND VPWR heichips25_can_lehmann_fsm/net991
+ heichips25_can_lehmann_fsm__3019_/Q clknet_leaf_21_clk sg13g2_dfrbpq_1
Xheichips25_sap3__2350_ heichips25_sap3/_1771_ net10 heichips25_sap3/_1770_ VPWR VGND
+ sg13g2_nand2_1
XFILLER_28_641 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2281_ heichips25_sap3/_1702_ heichips25_sap3/net270 heichips25_sap3/_1617_
+ VPWR VGND sg13g2_nand2_1
XFILLER_15_302 VPWR VGND sg13g2_fill_2
XFILLER_43_622 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__4020_ heichips25_sap3/net446 VGND VPWR heichips25_sap3/_0161_ heichips25_sap3__4020_/Q
+ clkload19/A sg13g2_dfrbpq_1
XFILLER_15_357 VPWR VGND sg13g2_decap_8
XFILLER_15_368 VPWR VGND sg13g2_fill_1
XFILLER_16_869 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3804_ VGND VPWR heichips25_sap3__4007_/Q heichips25_sap3/_1278_
+ heichips25_sap3/_1312_ heichips25_sap3/net291 sg13g2_a21oi_1
Xheichips25_sap3__1996_ VPWR heichips25_sap3/_1422_ heichips25_sap3__4002_/Q VGND
+ sg13g2_inv_1
Xheichips25_sap3__3735_ heichips25_sap3__4029_/Q heichips25_sap3__4033_/Q heichips25_sap3__4034_/Q
+ heichips25_sap3__4035_/Q heichips25_sap3__4036_/Q heichips25_sap3__4030_/Q heichips25_sap3/_1252_
+ VPWR VGND sg13g2_mux4_1
Xheichips25_sap3__3666_ VPWR VGND heichips25_sap3/_0888_ heichips25_sap3/_1209_ heichips25_sap3/_1210_
+ heichips25_sap3/net96 heichips25_sap3/_1211_ heichips25_sap3/_0971_ sg13g2_a221oi_1
Xheichips25_sap3__2617_ heichips25_sap3/_0287_ heichips25_sap3/net1064 heichips25_sap3/_1433_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__3597_ heichips25_sap3/_0111_ heichips25_sap3/_1130_ heichips25_sap3/_1170_
+ heichips25_sap3/net101 heichips25_sap3/_1424_ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2548_ heichips25_sap3/_0223_ VPWR heichips25_sap3/_0224_ VGND heichips25_sap3/_1802_
+ uio_out_sap3\[0\] sg13g2_o21ai_1
Xheichips25_sap3__2479_ heichips25_sap3/_1884_ heichips25_sap3/net168 heichips25_sap3/_1892_
+ VPWR VGND sg13g2_nor2b_1
XFILLER_18_195 VPWR VGND sg13g2_fill_2
XFILLER_34_677 VPWR VGND sg13g2_fill_1
XFILLER_33_121 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2321_ VGND VPWR heichips25_can_lehmann_fsm/_0971_ heichips25_can_lehmann_fsm/net363
+ heichips25_can_lehmann_fsm/_0060_ heichips25_can_lehmann_fsm/_0626_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2252_ VGND VPWR heichips25_can_lehmann_fsm/net898 heichips25_can_lehmann_fsm/net170
+ heichips25_can_lehmann_fsm/_0572_ heichips25_can_lehmann_fsm/_0571_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2183_ heichips25_can_lehmann_fsm/net325 VPWR heichips25_can_lehmann_fsm/_0518_
+ VGND heichips25_can_lehmann_fsm/net1236 heichips25_can_lehmann_fsm/net160 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2858__780 VPWR VGND net779 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2889__718 VPWR VGND net717 sg13g2_tiehi
XFILLER_5_1028 VPWR VGND sg13g2_fill_1
XFILLER_5_1017 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1967_ heichips25_can_lehmann_fsm/_0327_ heichips25_can_lehmann_fsm__2781_/Q
+ heichips25_can_lehmann_fsm/_1065_ VPWR VGND sg13g2_xnor2_1
Xheichips25_sap3_hold1122 heichips25_sap3__4050_/Q VPWR VGND heichips25_sap3/net1121
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__1898_ heichips25_can_lehmann_fsm/_1209_ heichips25_can_lehmann_fsm/_1210_
+ heichips25_can_lehmann_fsm/_1208_ heichips25_can_lehmann_fsm/_1211_ VPWR VGND sg13g2_nand3_1
Xheichips25_sap3_hold1144 heichips25_sap3__4053_/Q VPWR VGND heichips25_sap3/net1143
+ sg13g2_dlygate4sd3_1
XFILLER_24_176 VPWR VGND sg13g2_fill_1
Xheichips25_sap3_hold1177 heichips25_sap3__4029_/Q VPWR VGND heichips25_sap3/net1176
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__2519_ VGND VPWR heichips25_can_lehmann_fsm/_0918_ heichips25_can_lehmann_fsm/net417
+ heichips25_can_lehmann_fsm/_0159_ heichips25_can_lehmann_fsm/_0725_ sg13g2_a21oi_1
XFILLER_21_21 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm_fanout492 heichips25_can_lehmann_fsm/net493 heichips25_can_lehmann_fsm/net492
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout470 heichips25_can_lehmann_fsm/net503 heichips25_can_lehmann_fsm/net470
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout481 heichips25_can_lehmann_fsm/net490 heichips25_can_lehmann_fsm/net481
+ VPWR VGND sg13g2_buf_1
Xheichips25_sap3__3520_ heichips25_sap3/_1112_ VPWR heichips25_sap3/_1113_ VGND net46
+ heichips25_sap3/_1087_ sg13g2_o21ai_1
XFILLER_0_787 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3451_ uio_out_sap3\[0\] heichips25_sap3/_1053_ heichips25_sap3/_1055_
+ heichips25_sap3/_1056_ VPWR VGND sg13g2_or3_1
Xheichips25_sap3__3382_ heichips25_sap3/_0986_ heichips25_sap3/_0987_ heichips25_sap3/_0988_
+ heichips25_sap3/_0989_ heichips25_sap3/_0990_ VPWR VGND sg13g2_and4_1
Xheichips25_sap3__2402_ heichips25_sap3/_1817_ heichips25_sap3/_1819_ heichips25_sap3/_1742_
+ heichips25_sap3/_1821_ VPWR VGND heichips25_sap3/_1820_ sg13g2_nand4_1
Xheichips25_sap3__2333_ heichips25_sap3/net244 heichips25_sap3/_1530_ heichips25_sap3/_1531_
+ heichips25_sap3/_1754_ VPWR VGND sg13g2_nor3_1
XFILLER_44_931 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2264_ heichips25_sap3/_1503_ heichips25_sap3/net242 heichips25_sap3/_1522_
+ heichips25_sap3/_1526_ heichips25_sap3/_1685_ VPWR VGND sg13g2_nor4_1
XFILLER_28_493 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__4003_ heichips25_sap3/net456 VGND VPWR heichips25_sap3/_0144_ heichips25_sap3__4003_/Q
+ heichips25_sap3__4003_/CLK sg13g2_dfrbpq_1
Xheichips25_sap3__2195_ heichips25_sap3/_1616_ heichips25_sap3/net237 heichips25_sap3/_1613_
+ VPWR VGND sg13g2_nand2_1
XFILLER_31_669 VPWR VGND sg13g2_fill_2
XFILLER_12_883 VPWR VGND sg13g2_fill_1
XFILLER_11_371 VPWR VGND sg13g2_fill_1
XFILLER_7_386 VPWR VGND sg13g2_fill_2
X_24__510 VPWR VGND net509 sg13g2_tielo
Xheichips25_sap3__1979_ VPWR heichips25_sap3/_1405_ heichips25_sap3__4016_/Q VGND
+ sg13g2_inv_1
Xheichips25_sap3__3718_ heichips25_sap3/_1242_ VPWR heichips25_sap3/_0160_ VGND heichips25_sap3/_1393_
+ heichips25_sap3/net117 sg13g2_o21ai_1
XFILLER_30_4 VPWR VGND sg13g2_fill_1
XFILLER_39_725 VPWR VGND sg13g2_fill_2
XFILLER_38_202 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3649_ VPWR VGND heichips25_sap3/_1197_ heichips25_sap3/net112 heichips25_sap3/_1196_
+ heichips25_sap3/net98 heichips25_sap3/_1198_ heichips25_sap3/_0875_ sg13g2_a221oi_1
XFILLER_16_2 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2870_ net755 VGND VPWR heichips25_can_lehmann_fsm/_0095_
+ heichips25_can_lehmann_fsm__2870_/Q clknet_leaf_20_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1821_ VPWR VGND heichips25_can_lehmann_fsm/_1114_ heichips25_can_lehmann_fsm/_1131_
+ heichips25_can_lehmann_fsm/_1135_ heichips25_can_lehmann_fsm/_1075_ heichips25_can_lehmann_fsm/_1137_
+ heichips25_can_lehmann_fsm/_1134_ sg13g2_a221oi_1
XFILLER_47_780 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1752_ heichips25_can_lehmann_fsm__2789_/Q heichips25_can_lehmann_fsm__2788_/Q
+ heichips25_can_lehmann_fsm/_1068_ heichips25_can_lehmann_fsm/_1069_ heichips25_can_lehmann_fsm/_1072_
+ VPWR VGND sg13g2_or4_1
Xheichips25_can_lehmann_fsm__1683_ heichips25_can_lehmann_fsm/_1007_ heichips25_can_lehmann_fsm/net331
+ heichips25_can_lehmann_fsm__3041_/Q heichips25_can_lehmann_fsm/net313 heichips25_can_lehmann_fsm__2921_/Q
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2304_ VGND VPWR heichips25_can_lehmann_fsm/net1085 heichips25_can_lehmann_fsm/net173
+ heichips25_can_lehmann_fsm/_0614_ heichips25_can_lehmann_fsm/_0613_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2235_ heichips25_can_lehmann_fsm/net1212 heichips25_can_lehmann_fsm/net170
+ heichips25_can_lehmann_fsm/_0558_ VPWR VGND sg13g2_nor2_1
Xheichips25_can_lehmann_fsm__2166_ VPWR VGND net12 heichips25_can_lehmann_fsm/_0497_
+ heichips25_can_lehmann_fsm/_0499_ heichips25_can_lehmann_fsm/net1093 heichips25_can_lehmann_fsm/_0504_
+ heichips25_can_lehmann_fsm/net175 sg13g2_a221oi_1
Xheichips25_can_lehmann_fsm__2097_ VPWR VGND heichips25_can_lehmann_fsm/_0437_ heichips25_can_lehmann_fsm/net183
+ heichips25_can_lehmann_fsm/net186 heichips25_can_lehmann_fsm/net1268 heichips25_can_lehmann_fsm/_0438_
+ heichips25_can_lehmann_fsm/_0307_ sg13g2_a221oi_1
XFILLER_17_408 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2999_ net601 VGND VPWR heichips25_can_lehmann_fsm/_0224_
+ heichips25_can_lehmann_fsm__2999_/Q clknet_leaf_6_clk sg13g2_dfrbpq_1
Xheichips25_sap3_fanout341 heichips25_sap3/net1276 heichips25_sap3/net341 VPWR VGND
+ sg13g2_buf_1
XFILLER_16_43 VPWR VGND sg13g2_decap_4
XFILLER_25_452 VPWR VGND sg13g2_decap_4
XFILLER_26_964 VPWR VGND sg13g2_fill_2
XFILLER_12_102 VPWR VGND sg13g2_decap_8
XFILLER_12_124 VPWR VGND sg13g2_decap_8
XFILLER_40_477 VPWR VGND sg13g2_decap_8
XFILLER_40_455 VPWR VGND sg13g2_fill_1
XFILLER_8_117 VPWR VGND sg13g2_decap_4
XFILLER_8_106 VPWR VGND sg13g2_decap_4
XFILLER_32_31 VPWR VGND sg13g2_decap_8
XFILLER_8_139 VPWR VGND sg13g2_fill_2
XFILLER_8_128 VPWR VGND sg13g2_fill_1
XFILLER_32_42 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2951_ heichips25_sap3/_0588_ heichips25_sap3/_0563_ heichips25_sap3/_0589_
+ VPWR VGND sg13g2_xor2_1
XFILLER_4_323 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2882_ heichips25_sap3/_0522_ heichips25_sap3/_0379_ heichips25_sap3/_0523_
+ VPWR VGND sg13g2_xor2_1
Xheichips25_sap3__3503_ heichips25_sap3/net106 heichips25_sap3/_1098_ heichips25_sap3/_1099_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__3434_ VPWR heichips25_sap3/_1040_ heichips25_sap3/_1039_ VGND sg13g2_inv_1
XFILLER_36_717 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3365_ heichips25_sap3/net96 VPWR heichips25_sap3/_0974_ VGND heichips25_sap3/net124
+ heichips25_sap3/_0973_ sg13g2_o21ai_1
XFILLER_35_249 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2316_ heichips25_sap3/_1695_ heichips25_sap3/_1736_ heichips25_sap3/_1737_
+ VPWR VGND sg13g2_and2_1
Xheichips25_sap3__3296_ VPWR VGND heichips25_sap3/_0907_ heichips25_sap3/_0732_ heichips25_sap3/_0906_
+ heichips25_sap3/net122 heichips25_sap3/_0908_ heichips25_sap3/_0905_ sg13g2_a221oi_1
XFILLER_32_901 VPWR VGND sg13g2_fill_1
XFILLER_44_772 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2247_ VGND VPWR heichips25_sap3/net266 heichips25_sap3/net262 heichips25_sap3/_1668_
+ heichips25_sap3/_1365_ sg13g2_a21oi_1
XFILLER_43_293 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2178_ heichips25_sap3/_1519_ heichips25_sap3/net225 heichips25_sap3/_1599_
+ VPWR VGND sg13g2_nor2_1
XFILLER_12_680 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2020_ VGND VPWR heichips25_can_lehmann_fsm/_0369_ heichips25_can_lehmann_fsm/_0371_
+ heichips25_can_lehmann_fsm/_0013_ heichips25_can_lehmann_fsm/_0372_ sg13g2_a21oi_1
XFILLER_4_890 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2922_ net647 VGND VPWR heichips25_can_lehmann_fsm/_0147_
+ heichips25_can_lehmann_fsm__2922_/Q clknet_leaf_21_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2853_ net789 VGND VPWR heichips25_can_lehmann_fsm/_0078_
+ heichips25_can_lehmann_fsm__2853_/Q clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_39_588 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__1804_ heichips25_can_lehmann_fsm/net338 heichips25_can_lehmann_fsm/_0992_
+ heichips25_can_lehmann_fsm__2924_/Q heichips25_can_lehmann_fsm/_1120_ VPWR VGND
+ sg13g2_nand3_1
XFILLER_26_216 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2784_ net638 VGND VPWR heichips25_can_lehmann_fsm/net1235
+ heichips25_can_lehmann_fsm__2784_/Q clknet_leaf_5_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1735_ heichips25_can_lehmann_fsm/_1055_ VPWR uo_out_fsm\[3\]
+ VGND heichips25_can_lehmann_fsm/_1030_ heichips25_can_lehmann_fsm/_1054_ sg13g2_o21ai_1
XFILLER_23_934 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1666_ heichips25_can_lehmann_fsm/net350 heichips25_can_lehmann_fsm/_0989_
+ heichips25_can_lehmann_fsm/_0990_ VPWR VGND sg13g2_and2_1
XFILLER_34_271 VPWR VGND sg13g2_decap_8
XFILLER_34_293 VPWR VGND sg13g2_decap_8
XFILLER_10_606 VPWR VGND sg13g2_decap_8
XFILLER_23_978 VPWR VGND sg13g2_fill_1
XFILLER_22_488 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1597_ VPWR heichips25_can_lehmann_fsm/_0921_ heichips25_can_lehmann_fsm/net1062
+ VGND sg13g2_inv_1
XFILLER_5_109 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2218_ heichips25_can_lehmann_fsm/_0545_ heichips25_can_lehmann_fsm/net165
+ heichips25_can_lehmann_fsm/_0544_ heichips25_can_lehmann_fsm/net176 heichips25_can_lehmann_fsm/net1034
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2149_ heichips25_can_lehmann_fsm/_0488_ heichips25_can_lehmann_fsm/_0484_
+ heichips25_can_lehmann_fsm/_0487_ heichips25_can_lehmann_fsm/net301 heichips25_can_lehmann_fsm/_0948_
+ VPWR VGND sg13g2_a22oi_1
XFILLER_49_308 VPWR VGND sg13g2_decap_4
XFILLER_17_249 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3150_ heichips25_sap3/net152 heichips25_sap3/_0762_ heichips25_sap3/_0763_
+ VPWR VGND sg13g2_and2_1
Xheichips25_sap3__2101_ heichips25_sap3/net267 heichips25_sap3/_1438_ heichips25_sap3/_1488_
+ heichips25_sap3/_1522_ VGND VPWR heichips25_sap3/_1511_ sg13g2_nor4_2
Xheichips25_sap3__3081_ VGND VPWR heichips25_sap3/net220 heichips25_sap3/_0689_ heichips25_sap3/_0694_
+ heichips25_sap3/net249 sg13g2_a21oi_1
Xheichips25_sap3__2032_ heichips25_sap3/_1444_ heichips25_sap3/_1450_ heichips25_sap3/_1453_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_can_lehmann_fsm_hold1250 heichips25_can_lehmann_fsm__2780_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1249 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__2943__564 VPWR VGND net563 sg13g2_tiehi
XFILLER_9_415 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm_hold1272 heichips25_can_lehmann_fsm/_0025_ VPWR VGND heichips25_can_lehmann_fsm/net1271
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1261 heichips25_can_lehmann_fsm__2781_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1260 sg13g2_dlygate4sd3_1
XFILLER_13_488 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3983_ heichips25_sap3/net439 VGND VPWR heichips25_sap3/_0124_ heichips25_sap3__3983_/Q
+ heichips25_sap3__4015_/CLK sg13g2_dfrbpq_1
XFILLER_5_610 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2934_ heichips25_sap3/_0571_ VPWR heichips25_sap3/_0573_ VGND heichips25_sap3/_0341_
+ heichips25_sap3/_0572_ sg13g2_o21ai_1
Xheichips25_sap3__2865_ heichips25_sap3/_0506_ VPWR heichips25_sap3/_0507_ VGND heichips25_sap3/_0502_
+ heichips25_sap3/_0505_ sg13g2_o21ai_1
XFILLER_4_175 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2796_ heichips25_sap3/_1881_ heichips25_sap3/_1884_ heichips25_sap3/_1880_
+ heichips25_sap3/_0441_ VPWR VGND heichips25_sap3/net168 sg13g2_nand4_1
XFILLER_4_46 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2915__666 VPWR VGND net665 sg13g2_tiehi
XFILLER_4_79 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3417_ heichips25_sap3/_1024_ heichips25_sap3/_0999_ heichips25_sap3/_1014_
+ VPWR VGND sg13g2_xnor2_1
Xheichips25_sap3__3348_ heichips25_sap3/net55 heichips25_sap3/_0954_ heichips25_sap3/_0956_
+ heichips25_sap3/_0958_ VPWR VGND sg13g2_nor3_1
XFILLER_16_260 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3279_ heichips25_sap3/_0891_ heichips25_sap3__3932_/Q heichips25_sap3/net55
+ VPWR VGND sg13g2_nand2_1
XFILLER_31_241 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2922__648 VPWR VGND net647 sg13g2_tiehi
XFILLER_8_470 VPWR VGND sg13g2_decap_8
XFILLER_8_481 VPWR VGND sg13g2_fill_1
XFILLER_8_492 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__3052_ net766 VGND VPWR heichips25_can_lehmann_fsm/net1156
+ heichips25_can_lehmann_fsm__3052_/Q clknet_leaf_11_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2003_ heichips25_can_lehmann_fsm/_0358_ heichips25_can_lehmann_fsm__2786_/Q
+ heichips25_can_lehmann_fsm/_1068_ VPWR VGND sg13g2_xnor2_1
Xheichips25_can_lehmann_fsm__2816__575 VPWR VGND net574 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2905_ net685 VGND VPWR heichips25_can_lehmann_fsm/net1042
+ heichips25_can_lehmann_fsm__2905_/Q clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_27_503 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2836_ net534 VGND VPWR heichips25_can_lehmann_fsm/_0061_
+ heichips25_can_lehmann_fsm__2836_/Q clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_27_558 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2767_ VGND VPWR heichips25_can_lehmann_fsm/_0853_ heichips25_can_lehmann_fsm/net412
+ heichips25_can_lehmann_fsm/_0283_ heichips25_can_lehmann_fsm/_0849_ sg13g2_a21oi_1
Xclkbuf_5_29__f_heichips25_sap3\_sap_3_inst.alu_inst.clk clkload28/A clknet_4_14_0_heichips25_sap3\/sap_3_inst.alu_inst.clk
+ VPWR VGND sg13g2_buf_16
Xheichips25_can_lehmann_fsm__1718_ heichips25_can_lehmann_fsm/_1040_ VPWR uo_out_fsm\[1\]
+ VGND heichips25_can_lehmann_fsm/_1010_ heichips25_can_lehmann_fsm/_1039_ sg13g2_o21ai_1
XFILLER_23_731 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2698_ heichips25_can_lehmann_fsm/net494 VPWR heichips25_can_lehmann_fsm/_0815_
+ VGND heichips25_can_lehmann_fsm/net1114 heichips25_can_lehmann_fsm/net382 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__1649_ VPWR heichips25_can_lehmann_fsm/_0973_ heichips25_can_lehmann_fsm/net1182
+ VGND sg13g2_inv_1
XFILLER_11_926 VPWR VGND sg13g2_fill_2
XFILLER_22_263 VPWR VGND sg13g2_decap_8
XFILLER_8_4 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2650_ heichips25_sap3/_0316_ VPWR heichips25_sap3/_0317_ VGND heichips25_sap3/_1875_
+ heichips25_sap3/_0314_ sg13g2_o21ai_1
XFILLER_49_116 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2581_ heichips25_sap3/_0254_ heichips25_sap3/net74 heichips25_sap3__3997_/Q
+ heichips25_sap3/net79 heichips25_sap3__4021_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_49_149 VPWR VGND sg13g2_fill_2
XFILLER_38_63 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3202_ heichips25_sap3/_0811_ heichips25_sap3/_0812_ heichips25_sap3/_0813_
+ heichips25_sap3/_0814_ heichips25_sap3/_0815_ VPWR VGND sg13g2_and4_1
XFILLER_45_366 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3133_ heichips25_sap3/_0746_ heichips25_sap3/_0662_ heichips25_sap3/_0745_
+ VPWR VGND sg13g2_nand2b_1
XFILLER_33_506 VPWR VGND sg13g2_decap_8
XFILLER_33_517 VPWR VGND sg13g2_fill_2
XFILLER_33_528 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3064_ heichips25_sap3/net258 heichips25_sap3/_1448_ heichips25_sap3/net226
+ heichips25_sap3/_1722_ heichips25_sap3/_0677_ VPWR VGND sg13g2_or4_1
XFILLER_13_230 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2015_ heichips25_sap3/net267 heichips25_sap3/net264 heichips25_sap3/_1436_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_can_lehmann_fsm_hold1080 heichips25_can_lehmann_fsm__2936_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1079 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1091 heichips25_can_lehmann_fsm__2996_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1090 sg13g2_dlygate4sd3_1
Xclkload15 clkload15/Y clknet_leaf_10_clk VPWR VGND sg13g2_inv_2
XFILLER_9_278 VPWR VGND sg13g2_fill_1
Xclkload26 VPWR clkload26/Y clkload26/A VGND sg13g2_inv_1
XFILLER_6_963 VPWR VGND sg13g2_fill_1
XFILLER_10_992 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3966_ heichips25_sap3/net438 VGND VPWR heichips25_sap3/_0107_ heichips25_sap3__3966_/Q
+ heichips25_sap3__4014_/CLK sg13g2_dfrbpq_1
XFILLER_6_996 VPWR VGND sg13g2_decap_4
XFILLER_5_462 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2917_ VGND VPWR heichips25_sap3/net65 heichips25_sap3/_0545_ heichips25_sap3/_0557_
+ heichips25_sap3/net203 sg13g2_a21oi_1
Xheichips25_sap3__3897_ heichips25_sap3/net449 VGND VPWR heichips25_sap3/_0038_ heichips25_sap3__3897_/Q
+ net821 sg13g2_dfrbpq_1
Xheichips25_sap3__2848_ heichips25_sap3/_0491_ heichips25_sap3/_0490_ heichips25_sap3/_0340_
+ heichips25_sap3/_0489_ heichips25_sap3/_0338_ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2779_ heichips25_sap3/_0336_ VPWR heichips25_sap3/_0039_ VGND heichips25_sap3/_0423_
+ heichips25_sap3/_0424_ sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2621_ VGND VPWR heichips25_can_lehmann_fsm/_0892_ heichips25_can_lehmann_fsm/net375
+ heichips25_can_lehmann_fsm/_0210_ heichips25_can_lehmann_fsm/_0776_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2552_ heichips25_can_lehmann_fsm/net472 VPWR heichips25_can_lehmann_fsm/_0742_
+ VGND heichips25_can_lehmann_fsm__2950_/Q heichips25_can_lehmann_fsm/net365 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2483_ VGND VPWR heichips25_can_lehmann_fsm/_0927_ heichips25_can_lehmann_fsm/net409
+ heichips25_can_lehmann_fsm/_0141_ heichips25_can_lehmann_fsm/_0707_ sg13g2_a21oi_1
Xclkload9 VPWR clkload9/Y clknet_leaf_15_clk VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__3057__558 VPWR VGND net557 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__3035_ net549 VGND VPWR heichips25_can_lehmann_fsm/_0260_
+ heichips25_can_lehmann_fsm__3035_/Q clknet_leaf_18_clk sg13g2_dfrbpq_1
XFILLER_28_834 VPWR VGND sg13g2_decap_4
XFILLER_42_303 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2868__760 VPWR VGND net759 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2819_ net568 VGND VPWR heichips25_can_lehmann_fsm/net1175
+ heichips25_can_lehmann_fsm__2819_/Q clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_42_336 VPWR VGND sg13g2_decap_8
XFILLER_42_325 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm_hold900 heichips25_can_lehmann_fsm/_0079_ VPWR VGND heichips25_can_lehmann_fsm/net899
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold944 heichips25_can_lehmann_fsm/_0084_ VPWR VGND heichips25_can_lehmann_fsm/net943
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold922 heichips25_can_lehmann_fsm__2968_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net921 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold933 heichips25_can_lehmann_fsm/_0231_ VPWR VGND heichips25_can_lehmann_fsm/net932
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold911 heichips25_can_lehmann_fsm/_0135_ VPWR VGND heichips25_can_lehmann_fsm/net910
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold966 heichips25_can_lehmann_fsm__2857_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net965 sg13g2_dlygate4sd3_1
XFILLER_23_594 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_hold977 heichips25_can_lehmann_fsm__2884_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net976 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold999 heichips25_can_lehmann_fsm__3017_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net998 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold988 heichips25_can_lehmann_fsm__2869_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net987 sg13g2_dlygate4sd3_1
Xheichips25_sap3__3820_ heichips25_sap3/net340 heichips25_sap3/net1011 heichips25_sap3/_1326_
+ heichips25_sap3/_0178_ VPWR VGND sg13g2_a21o_1
Xheichips25_sap3__3751_ heichips25_sap3/_1263_ heichips25_sap3/net293 heichips25_sap3__3987_/Q
+ heichips25_sap3/_1259_ heichips25_sap3__3979_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_3_944 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2702_ heichips25_sap3/_0348_ heichips25_sap3/net274 heichips25_sap3__3922_/Q
+ VPWR VGND sg13g2_nand2_1
XFILLER_2_410 VPWR VGND sg13g2_fill_2
XFILLER_46_1021 VPWR VGND sg13g2_decap_8
XFILLER_3_977 VPWR VGND sg13g2_decap_8
XFILLER_2_443 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3682_ VGND VPWR heichips25_sap3/net60 heichips25_sap3/net99 heichips25_sap3/_1223_
+ heichips25_sap3/net113 sg13g2_a21oi_1
Xheichips25_sap3__2633_ heichips25_sap3/_1718_ heichips25_sap3/_1774_ heichips25_sap3/_1573_
+ heichips25_sap3/_0300_ VPWR VGND heichips25_sap3/_0299_ sg13g2_nand4_1
XFILLER_49_95 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2564_ heichips25_sap3/_0239_ heichips25_sap3/net85 heichips25_sap3__3958_/Q
+ heichips25_sap3/net88 heichips25_sap3__3950_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_19_801 VPWR VGND sg13g2_fill_2
XFILLER_19_867 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2495_ VPWR VGND heichips25_sap3/_1907_ heichips25_sap3/_1654_ heichips25_sap3/_1904_
+ heichips25_sap3/_1385_ heichips25_sap3/_1908_ heichips25_sap3/net89 sg13g2_a221oi_1
XFILLER_18_377 VPWR VGND sg13g2_fill_1
XFILLER_34_859 VPWR VGND sg13g2_fill_2
XFILLER_33_325 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3116_ heichips25_sap3/_0723_ heichips25_sap3/_0724_ heichips25_sap3/_0728_
+ heichips25_sap3/_0729_ VPWR VGND sg13g2_nor3_1
Xheichips25_sap3__3047_ heichips25_sap3/_0660_ heichips25_sap3/_1364_ heichips25_sap3/_1451_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__3949_ heichips25_sap3/net433 VGND VPWR heichips25_sap3/_0090_ heichips25_sap3__3949_/Q
+ heichips25_sap3__4013_/CLK sg13g2_dfrbpq_1
XFILLER_5_292 VPWR VGND sg13g2_fill_2
Xinput2 rst_n net2 VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm__1983_ heichips25_can_lehmann_fsm/net185 VPWR heichips25_can_lehmann_fsm/_0341_
+ VGND heichips25_can_lehmann_fsm/_0339_ heichips25_can_lehmann_fsm/_0340_ sg13g2_o21ai_1
XFILLER_28_108 VPWR VGND sg13g2_fill_2
XFILLER_37_686 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2604_ heichips25_can_lehmann_fsm/net491 VPWR heichips25_can_lehmann_fsm/_0768_
+ VGND heichips25_can_lehmann_fsm/net930 heichips25_can_lehmann_fsm/net380 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2535_ VGND VPWR heichips25_can_lehmann_fsm/_0914_ heichips25_can_lehmann_fsm/net395
+ heichips25_can_lehmann_fsm/_0167_ heichips25_can_lehmann_fsm/_0733_ sg13g2_a21oi_1
XFILLER_20_531 VPWR VGND sg13g2_fill_2
XFILLER_32_391 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2466_ heichips25_can_lehmann_fsm/net498 VPWR heichips25_can_lehmann_fsm/_0699_
+ VGND heichips25_can_lehmann_fsm/net903 heichips25_can_lehmann_fsm/net426 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2397_ VGND VPWR heichips25_can_lehmann_fsm/_0952_ heichips25_can_lehmann_fsm/net390
+ heichips25_can_lehmann_fsm/_0098_ heichips25_can_lehmann_fsm/_0664_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__3018_ net738 VGND VPWR heichips25_can_lehmann_fsm/_0243_
+ heichips25_can_lehmann_fsm__3018_/Q clknet_leaf_20_clk sg13g2_dfrbpq_1
XFILLER_0_936 VPWR VGND sg13g2_decap_8
XFILLER_48_918 VPWR VGND sg13g2_fill_1
XFILLER_19_10 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2280_ heichips25_sap3/_1701_ heichips25_sap3/_1700_ heichips25_sap3/_1564_
+ heichips25_sap3/_1696_ heichips25_sap3/_1539_ VPWR VGND sg13g2_a22oi_1
XFILLER_27_152 VPWR VGND sg13g2_fill_2
XFILLER_35_42 VPWR VGND sg13g2_fill_2
XFILLER_15_314 VPWR VGND sg13g2_decap_8
XFILLER_27_185 VPWR VGND sg13g2_decap_8
XFILLER_42_155 VPWR VGND sg13g2_decap_8
XFILLER_7_535 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3803_ heichips25_sap3/_1311_ heichips25_sap3/_1282_ heichips25_sap3__3951_/Q
+ heichips25_sap3/_1270_ heichips25_sap3__4023_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__1995_ VPWR heichips25_sap3/_1421_ heichips25_sap3__4018_/Q VGND
+ sg13g2_inv_1
Xheichips25_sap3__3734_ VGND VPWR heichips25_sap3/_1248_ heichips25_sap3/_1250_ heichips25_sap3/_1251_
+ heichips25_sap3/_1432_ sg13g2_a21oi_1
Xheichips25_sap3__3665_ heichips25_sap3/_0969_ VPWR heichips25_sap3/_1210_ VGND heichips25_sap3/_0945_
+ heichips25_sap3/_0965_ sg13g2_o21ai_1
Xheichips25_sap3__2616_ heichips25_sap3/_1359_ heichips25_sap3/net1019 heichips25_sap3/_0286_
+ VPWR VGND sg13g2_nor2_1
XFILLER_2_284 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3596_ heichips25_sap3/net101 heichips25_sap3/_1131_ heichips25_sap3/_1169_
+ heichips25_sap3/_1170_ VPWR VGND sg13g2_nor3_1
Xheichips25_sap3__2547_ heichips25_sap3/_1717_ heichips25_sap3/_1878_ heichips25_sap3/_0222_
+ heichips25_sap3/_0223_ VPWR VGND sg13g2_nor3_1
Xheichips25_sap3__2478_ heichips25_sap3/_1890_ VPWR heichips25_sap3/_1891_ VGND heichips25_sap3/_1518_
+ heichips25_sap3/_1560_ sg13g2_o21ai_1
XFILLER_34_623 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2320_ heichips25_can_lehmann_fsm/net474 VPWR heichips25_can_lehmann_fsm/_0626_
+ VGND heichips25_can_lehmann_fsm__2834_/Q heichips25_can_lehmann_fsm/net363 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2251_ VGND VPWR heichips25_can_lehmann_fsm/_1044_ heichips25_can_lehmann_fsm/_0570_
+ heichips25_can_lehmann_fsm/_0571_ heichips25_can_lehmann_fsm/net170 sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2182_ VPWR VGND net15 heichips25_can_lehmann_fsm/_0497_
+ heichips25_can_lehmann_fsm/_0499_ heichips25_can_lehmann_fsm/net933 heichips25_can_lehmann_fsm/_0517_
+ heichips25_can_lehmann_fsm/net175 sg13g2_a221oi_1
Xheichips25_can_lehmann_fsm__1966_ heichips25_can_lehmann_fsm__2781_/Q heichips25_can_lehmann_fsm/_1065_
+ heichips25_can_lehmann_fsm/_0326_ VPWR VGND sg13g2_nor2_1
Xheichips25_can_lehmann_fsm__1897_ heichips25_can_lehmann_fsm/_1210_ heichips25_can_lehmann_fsm/net314
+ heichips25_can_lehmann_fsm__2929_/Q heichips25_can_lehmann_fsm/net318 heichips25_can_lehmann_fsm__3001_/Q
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3_hold1145 heichips25_sap3/_0194_ VPWR VGND heichips25_sap3/net1144
+ sg13g2_dlygate4sd3_1
XFILLER_12_317 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2518_ heichips25_can_lehmann_fsm/net485 VPWR heichips25_can_lehmann_fsm/_0725_
+ VGND heichips25_can_lehmann_fsm__2934_/Q heichips25_can_lehmann_fsm/net417 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2449_ VGND VPWR heichips25_can_lehmann_fsm/_0935_ heichips25_can_lehmann_fsm/net359
+ heichips25_can_lehmann_fsm/_0124_ heichips25_can_lehmann_fsm/_0690_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2939__580 VPWR VGND net579 sg13g2_tiehi
Xheichips25_can_lehmann_fsm_fanout471 heichips25_can_lehmann_fsm/net475 heichips25_can_lehmann_fsm/net471
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout493 heichips25_can_lehmann_fsm/net496 heichips25_can_lehmann_fsm/net493
+ VPWR VGND sg13g2_buf_1
XFILLER_0_700 VPWR VGND sg13g2_decap_8
XFILLER_0_711 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm_fanout482 heichips25_can_lehmann_fsm/net484 heichips25_can_lehmann_fsm/net482
+ VPWR VGND sg13g2_buf_1
XFILLER_0_755 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3450_ VGND VPWR heichips25_sap3/_0736_ heichips25_sap3/net62 heichips25_sap3/_1055_
+ heichips25_sap3/_0731_ sg13g2_a21oi_1
Xheichips25_sap3__2401_ heichips25_sap3/_1820_ heichips25_sap3/net72 heichips25_sap3__3985_/Q
+ heichips25_sap3/net216 heichips25_sap3__4017_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3381_ heichips25_sap3/_0989_ heichips25_sap3/net104 heichips25_sap3__3944_/Q
+ heichips25_sap3/_0760_ heichips25_sap3__3960_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2332_ VGND VPWR heichips25_sap3/net249 heichips25_sap3/net225 heichips25_sap3/_1753_
+ heichips25_sap3/_1455_ sg13g2_a21oi_1
XFILLER_29_962 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2263_ heichips25_sap3/_1684_ heichips25_sap3/_1683_ heichips25_sap3/_1531_
+ heichips25_sap3/_1545_ heichips25_sap3/_1530_ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__4002_ heichips25_sap3/net442 VGND VPWR heichips25_sap3/_0143_ heichips25_sap3__4002_/Q
+ heichips25_sap3__4018_/CLK sg13g2_dfrbpq_1
XFILLER_44_954 VPWR VGND sg13g2_decap_4
XFILLER_15_111 VPWR VGND sg13g2_decap_8
XFILLER_15_122 VPWR VGND sg13g2_fill_2
XFILLER_15_144 VPWR VGND sg13g2_decap_8
XFILLER_43_475 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2194_ heichips25_sap3/_1615_ heichips25_sap3/net259 heichips25_sap3__3929_/Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_31_659 VPWR VGND sg13g2_fill_2
XFILLER_8_855 VPWR VGND sg13g2_fill_2
XFILLER_7_79 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__1978_ VPWR heichips25_sap3/_1404_ heichips25_sap3__3936_/Q VGND
+ sg13g2_inv_1
Xheichips25_sap3__3717_ heichips25_sap3/_1056_ heichips25_sap3/_1057_ heichips25_sap3/net117
+ heichips25_sap3/_1242_ VPWR VGND sg13g2_nand3_1
Xclkbuf_0_heichips25_sap3\_sap_3_inst.alu_inst.clk clknet_0_heichips25_sap3\/sap_3_inst.alu_inst.clk
+ heichips25_sap3/sap_3_inst.alu_inst.clk VPWR VGND sg13g2_buf_16
Xheichips25_sap3__3648_ uio_oe_sap3\[0\] heichips25_sap3/net98 heichips25_sap3/_1053_
+ heichips25_sap3/_1197_ VPWR VGND sg13g2_nor3_1
Xheichips25_sap3__3579_ VGND VPWR heichips25_sap3/net45 heichips25_sap3/net95 heichips25_sap3/_1157_
+ heichips25_sap3/_1156_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__1820_ heichips25_can_lehmann_fsm/_1136_ heichips25_can_lehmann_fsm/_1054_
+ heichips25_can_lehmann_fsm/_1123_ VPWR VGND sg13g2_nand2_1
Xheichips25_can_lehmann_fsm__1751_ heichips25_can_lehmann_fsm__2789_/Q heichips25_can_lehmann_fsm__2788_/Q
+ heichips25_can_lehmann_fsm/_1068_ heichips25_can_lehmann_fsm/_1069_ heichips25_can_lehmann_fsm/_1071_
+ VPWR VGND sg13g2_nor4_1
Xheichips25_can_lehmann_fsm__1682_ heichips25_can_lehmann_fsm/_1006_ heichips25_can_lehmann_fsm/net294
+ heichips25_can_lehmann_fsm__2969_/Q heichips25_can_lehmann_fsm/net310 heichips25_can_lehmann_fsm__3017_/Q
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2780__647 VPWR VGND net646 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2303_ heichips25_can_lehmann_fsm/net173 heichips25_can_lehmann_fsm/_0612_
+ heichips25_can_lehmann_fsm/_0613_ VPWR VGND sg13g2_nor2_1
Xheichips25_can_lehmann_fsm__2234_ heichips25_can_lehmann_fsm/_0557_ heichips25_can_lehmann_fsm/_0492_
+ heichips25_can_lehmann_fsm/_0461_ VPWR VGND sg13g2_nand2b_1
Xheichips25_can_lehmann_fsm__2165_ heichips25_can_lehmann_fsm/_0503_ heichips25_can_lehmann_fsm/net164
+ heichips25_can_lehmann_fsm/_0502_ VPWR VGND sg13g2_nand2_1
Xheichips25_can_lehmann_fsm__2096_ heichips25_can_lehmann_fsm/_0437_ heichips25_can_lehmann_fsm/net344
+ heichips25_can_lehmann_fsm/_1058_ VPWR VGND sg13g2_xnor2_1
XFILLER_29_258 VPWR VGND sg13g2_fill_2
XFILLER_29_269 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2998_ net609 VGND VPWR heichips25_can_lehmann_fsm/net856
+ heichips25_can_lehmann_fsm__2998_/Q clknet_leaf_6_clk sg13g2_dfrbpq_1
Xheichips25_sap3_fanout342 heichips25_sap3/net1071 heichips25_sap3/net342 VPWR VGND
+ sg13g2_buf_1
XFILLER_26_954 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1949_ heichips25_can_lehmann_fsm/_1215_ heichips25_can_lehmann_fsm/_1234_
+ heichips25_can_lehmann_fsm/_0312_ VPWR VGND sg13g2_nor2_1
XFILLER_41_935 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2826__555 VPWR VGND net554 sg13g2_tiehi
XFILLER_12_169 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2950_ heichips25_sap3/_0381_ heichips25_sap3/_0370_ heichips25_sap3/_0588_
+ VPWR VGND sg13g2_xor2_1
XFILLER_20_191 VPWR VGND sg13g2_decap_8
XFILLER_32_76 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2881_ heichips25_sap3/_0522_ heichips25_sap3/_0356_ heichips25_sap3/_0367_
+ VPWR VGND sg13g2_xnor2_1
XFILLER_5_869 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3502_ VGND VPWR heichips25_sap3/_0327_ heichips25_sap3/_1096_ heichips25_sap3/_1098_
+ heichips25_sap3/_1097_ sg13g2_a21oi_1
Xheichips25_sap3__3433_ heichips25_sap3/net96 VPWR heichips25_sap3/_1039_ VGND heichips25_sap3/net125
+ heichips25_sap3/_1038_ sg13g2_o21ai_1
XFILLER_48_567 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3364_ heichips25_sap3/_0872_ heichips25_sap3/_0972_ heichips25_sap3/_0973_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__2315_ VPWR VGND heichips25_sap3/_1730_ heichips25_sap3/_1711_ heichips25_sap3/_1715_
+ heichips25_sap3/_1708_ heichips25_sap3/_1736_ heichips25_sap3/_1707_ sg13g2_a221oi_1
XFILLER_44_740 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3295_ heichips25_sap3/_0907_ heichips25_sap3/_0327_ heichips25_sap3/net68
+ VPWR VGND sg13g2_nand2_1
XFILLER_44_762 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2246_ heichips25_sap3/_1601_ heichips25_sap3/net220 heichips25_sap3/_1667_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__2177_ heichips25_sap3/_1598_ heichips25_sap3/_1477_ heichips25_sap3/_1566_
+ VPWR VGND sg13g2_nand2_1
XFILLER_31_412 VPWR VGND sg13g2_fill_1
XFILLER_7_140 VPWR VGND sg13g2_decap_4
XFILLER_7_184 VPWR VGND sg13g2_decap_4
XFILLER_8_696 VPWR VGND sg13g2_decap_4
Xclkbuf_5_30__f_heichips25_sap3\_sap_3_inst.alu_inst.clk heichips25_sap3__3993_/CLK
+ clknet_4_15_0_heichips25_sap3\/sap_3_inst.alu_inst.clk VPWR VGND sg13g2_buf_16
Xheichips25_can_lehmann_fsm__2921_ net651 VGND VPWR heichips25_can_lehmann_fsm/net938
+ heichips25_can_lehmann_fsm__2921_/Q clknet_leaf_22_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2852_ net791 VGND VPWR heichips25_can_lehmann_fsm/net841
+ heichips25_can_lehmann_fsm__2852_/Q clknet_leaf_8_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1803_ heichips25_can_lehmann_fsm/_1119_ heichips25_can_lehmann_fsm__3044_/Q
+ heichips25_can_lehmann_fsm/net331 VPWR VGND sg13g2_nand2_1
Xheichips25_can_lehmann_fsm__2783_ net640 VGND VPWR heichips25_can_lehmann_fsm/_0008_
+ heichips25_can_lehmann_fsm__2783_/Q clknet_leaf_5_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1734_ heichips25_can_lehmann_fsm/_1055_ heichips25_can_lehmann_fsm/_1037_
+ heichips25_can_lehmann_fsm__2788_/Q heichips25_can_lehmann_fsm/_1032_ heichips25_can_lehmann_fsm__2797_/Q
+ VPWR VGND sg13g2_a22oi_1
XFILLER_22_412 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1665_ heichips25_can_lehmann_fsm/net351 heichips25_can_lehmann_fsm/net353
+ heichips25_can_lehmann_fsm/_0989_ VPWR VGND sg13g2_nor2b_1
Xheichips25_can_lehmann_fsm__1596_ VPWR heichips25_can_lehmann_fsm/_0920_ heichips25_can_lehmann_fsm/net858
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__2217_ heichips25_can_lehmann_fsm/_0544_ heichips25_can_lehmann_fsm/net1231
+ heichips25_can_lehmann_fsm/_1104_ VPWR VGND sg13g2_xnor2_1
XFILLER_1_316 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2148_ VPWR VGND heichips25_can_lehmann_fsm__2950_/Q heichips25_can_lehmann_fsm/_0486_
+ heichips25_can_lehmann_fsm/net306 heichips25_can_lehmann_fsm__3022_/Q heichips25_can_lehmann_fsm/_0487_
+ heichips25_can_lehmann_fsm/net312 sg13g2_a221oi_1
Xheichips25_can_lehmann_fsm__2079_ heichips25_can_lehmann_fsm/_1056_ VPWR heichips25_can_lehmann_fsm/_0423_
+ VGND heichips25_can_lehmann_fsm/_0976_ heichips25_can_lehmann_fsm/_0418_ sg13g2_o21ai_1
XFILLER_45_537 VPWR VGND sg13g2_fill_1
XFILLER_45_526 VPWR VGND sg13g2_fill_1
XFILLER_27_21 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2100_ heichips25_sap3/_1445_ heichips25_sap3/_1505_ heichips25_sap3/_1441_
+ heichips25_sap3/_1521_ VPWR VGND sg13g2_nand3_1
Xheichips25_sap3__3080_ heichips25_sap3/_0682_ heichips25_sap3/_0691_ heichips25_sap3/_0692_
+ heichips25_sap3/_0693_ VPWR VGND sg13g2_nor3_1
Xheichips25_sap3_fanout150 heichips25_sap3/_0751_ heichips25_sap3/net150 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3__2031_ heichips25_sap3/_1452_ heichips25_sap3/_1447_ heichips25_sap3/_1449_
+ VPWR VGND sg13g2_nand2_1
XFILLER_25_283 VPWR VGND sg13g2_fill_1
XFILLER_41_776 VPWR VGND sg13g2_fill_2
XFILLER_40_231 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm_hold1251 heichips25_can_lehmann_fsm/_0005_ VPWR VGND heichips25_can_lehmann_fsm/net1250
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1240 heichips25_can_lehmann_fsm/_0016_ VPWR VGND heichips25_can_lehmann_fsm/net1239
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1262 heichips25_can_lehmann_fsm/_0006_ VPWR VGND heichips25_can_lehmann_fsm/net1261
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1273 heichips25_can_lehmann_fsm__2868_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1272 sg13g2_dlygate4sd3_1
Xheichips25_sap3__3982_ heichips25_sap3/net439 VGND VPWR heichips25_sap3/_0123_ heichips25_sap3__3982_/Q
+ heichips25_sap3__4015_/CLK sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2878__740 VPWR VGND net739 sg13g2_tiehi
Xheichips25_sap3__2933_ heichips25_sap3/_0409_ heichips25_sap3/_0399_ heichips25_sap3/_0572_
+ VPWR VGND sg13g2_xor2_1
XFILLER_4_110 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2864_ VGND VPWR heichips25_sap3/_0502_ heichips25_sap3/_0505_ heichips25_sap3/_0506_
+ heichips25_sap3/_1869_ sg13g2_a21oi_1
Xheichips25_sap3__2795_ heichips25_sap3/_0440_ heichips25_sap3/_0439_ heichips25_sap3/_0437_
+ VPWR VGND sg13g2_nand2b_1
Xheichips25_can_lehmann_fsm__2950__536 VPWR VGND net535 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__3050__542 VPWR VGND net541 sg13g2_tiehi
XFILLER_49_843 VPWR VGND sg13g2_decap_8
XFILLER_0_360 VPWR VGND sg13g2_decap_8
XFILLER_0_371 VPWR VGND sg13g2_fill_2
XFILLER_49_865 VPWR VGND sg13g2_decap_8
XFILLER_49_854 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3416_ heichips25_sap3/_1022_ VPWR heichips25_sap3/_1023_ VGND heichips25_sap3/net123
+ heichips25_sap3/_1019_ sg13g2_o21ai_1
XFILLER_48_375 VPWR VGND sg13g2_fill_1
XFILLER_1_1010 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3347_ heichips25_sap3/_0957_ heichips25_sap3/_0819_ heichips25_sap3/_0854_
+ VPWR VGND sg13g2_xnor2_1
XFILLER_17_773 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3278_ heichips25_sap3/_0890_ VPWR heichips25_sap3/_0072_ VGND heichips25_sap3/_1392_
+ heichips25_sap3/_0747_ sg13g2_o21ai_1
Xheichips25_sap3__2229_ heichips25_sap3/_1473_ heichips25_sap3/_1648_ heichips25_sap3/_1649_
+ heichips25_sap3/_1650_ VPWR VGND sg13g2_nor3_1
XFILLER_31_220 VPWR VGND sg13g2_decap_8
XFILLER_31_264 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__3051_ net798 VGND VPWR heichips25_can_lehmann_fsm/_0276_
+ heichips25_can_lehmann_fsm__3051_/Q clknet_leaf_11_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2002_ VGND VPWR heichips25_can_lehmann_fsm/net1240 heichips25_can_lehmann_fsm/net188
+ heichips25_can_lehmann_fsm/_0357_ heichips25_can_lehmann_fsm/net191 sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2904_ net687 VGND VPWR heichips25_can_lehmann_fsm/net997
+ heichips25_can_lehmann_fsm__2904_/Q clknet_leaf_7_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2835_ net536 VGND VPWR heichips25_can_lehmann_fsm/net1094
+ heichips25_can_lehmann_fsm__2835_/Q clknet_leaf_5_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2766_ heichips25_can_lehmann_fsm/net485 VPWR heichips25_can_lehmann_fsm/_0849_
+ VGND heichips25_can_lehmann_fsm/net1148 heichips25_can_lehmann_fsm/net412 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__1717_ heichips25_can_lehmann_fsm/_1040_ heichips25_can_lehmann_fsm/_1037_
+ heichips25_can_lehmann_fsm__2786_/Q heichips25_can_lehmann_fsm/_1032_ heichips25_can_lehmann_fsm/net347
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2697_ VGND VPWR heichips25_can_lehmann_fsm/_0871_ heichips25_can_lehmann_fsm/net406
+ heichips25_can_lehmann_fsm/_0248_ heichips25_can_lehmann_fsm/_0814_ sg13g2_a21oi_1
Xfanout46 uio_out_sap3\[4\] net46 VPWR VGND sg13g2_buf_2
XFILLER_23_765 VPWR VGND sg13g2_decap_4
XFILLER_23_798 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__1648_ VPWR heichips25_can_lehmann_fsm/_0972_ net11 VGND
+ sg13g2_inv_1
Xheichips25_can_lehmann_fsm__1579_ VPWR heichips25_can_lehmann_fsm/_0903_ heichips25_can_lehmann_fsm/net1083
+ VGND sg13g2_inv_1
XFILLER_6_419 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2580_ VPWR VGND heichips25_sap3__3965_/Q heichips25_sap3/net89 heichips25_sap3/net82
+ heichips25_sap3__4005_/Q heichips25_sap3/_0253_ heichips25_sap3/net218 sg13g2_a221oi_1
XFILLER_38_42 VPWR VGND sg13g2_decap_8
XFILLER_45_312 VPWR VGND sg13g2_decap_8
XFILLER_45_345 VPWR VGND sg13g2_fill_2
XFILLER_45_323 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3201_ heichips25_sap3/_0814_ heichips25_sap3/net133 heichips25_sap3__3998_/Q
+ heichips25_sap3/net135 heichips25_sap3__3974_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3132_ VGND VPWR heichips25_sap3/_1454_ heichips25_sap3/_0744_ heichips25_sap3/_0745_
+ heichips25_sap3/net249 sg13g2_a21oi_1
Xheichips25_sap3__3063_ heichips25_sap3/net241 VPWR heichips25_sap3/_0676_ VGND heichips25_sap3/_0671_
+ heichips25_sap3/_0675_ sg13g2_o21ai_1
Xheichips25_sap3__2014_ VGND VPWR heichips25_sap3/_1435_ heichips25_sap3/net260 heichips25_sap3/net258
+ sg13g2_or2_1
Xheichips25_can_lehmann_fsm_hold1092 heichips25_can_lehmann_fsm__2964_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1091 sg13g2_dlygate4sd3_1
XFILLER_9_268 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm_hold1081 heichips25_can_lehmann_fsm__2873_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1080 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1070 heichips25_can_lehmann_fsm__2900_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1069 sg13g2_dlygate4sd3_1
Xclkload16 VPWR clkload16/Y clknet_leaf_11_clk VGND sg13g2_inv_1
XFILLER_10_960 VPWR VGND sg13g2_decap_8
XFILLER_10_971 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3965_ heichips25_sap3/net433 VGND VPWR heichips25_sap3/_0106_ heichips25_sap3__3965_/Q
+ heichips25_sap3__4013_/CLK sg13g2_dfrbpq_1
Xclkload27 VPWR clkload27/Y clkload27/A VGND sg13g2_inv_1
Xheichips25_sap3__2916_ heichips25_sap3/_0551_ VPWR heichips25_sap3/_0556_ VGND heichips25_sap3/_1869_
+ heichips25_sap3/_0555_ sg13g2_o21ai_1
Xheichips25_sap3__3896_ heichips25_sap3/net448 VGND VPWR heichips25_sap3/_0037_ heichips25_sap3__3896_/Q
+ net820 sg13g2_dfrbpq_1
Xheichips25_sap3__2847_ heichips25_sap3/_0490_ heichips25_sap3/_0402_ heichips25_sap3/_0403_
+ VPWR VGND sg13g2_xnor2_1
Xheichips25_sap3__2778_ heichips25_sap3/_0335_ VPWR heichips25_sap3/_0424_ VGND heichips25_sap3/_0345_
+ heichips25_sap3/_0371_ sg13g2_o21ai_1
Xheichips25_sap3__3875__820 VPWR net819 clkload27/A VGND sg13g2_inv_1
XFILLER_36_334 VPWR VGND sg13g2_fill_1
XFILLER_36_378 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2620_ heichips25_can_lehmann_fsm/net484 VPWR heichips25_can_lehmann_fsm/_0776_
+ VGND heichips25_can_lehmann_fsm/net984 heichips25_can_lehmann_fsm/net375 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2551_ VGND VPWR heichips25_can_lehmann_fsm/_0910_ heichips25_can_lehmann_fsm/net402
+ heichips25_can_lehmann_fsm/_0175_ heichips25_can_lehmann_fsm/_0741_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2482_ heichips25_can_lehmann_fsm/net482 VPWR heichips25_can_lehmann_fsm/_0707_
+ VGND heichips25_can_lehmann_fsm__2916_/Q heichips25_can_lehmann_fsm/net409 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__3034_ net565 VGND VPWR heichips25_can_lehmann_fsm/net1161
+ heichips25_can_lehmann_fsm__3034_/Q clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_39_150 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2818_ net570 VGND VPWR heichips25_can_lehmann_fsm/_0043_
+ heichips25_can_lehmann_fsm__2818_/Q clknet_leaf_8_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2749_ VGND VPWR heichips25_can_lehmann_fsm/_0857_ heichips25_can_lehmann_fsm/net381
+ heichips25_can_lehmann_fsm/_0274_ heichips25_can_lehmann_fsm/_0840_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm_hold901 heichips25_can_lehmann_fsm__2907_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net900 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold912 heichips25_can_lehmann_fsm__2852_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net911 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold934 heichips25_can_lehmann_fsm__2838_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net933 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold923 heichips25_can_lehmann_fsm__2867_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net922 sg13g2_dlygate4sd3_1
XFILLER_24_44 VPWR VGND sg13g2_decap_8
XFILLER_24_55 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_hold956 heichips25_can_lehmann_fsm__2891_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net955 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold945 heichips25_can_lehmann_fsm__3040_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net944 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold967 heichips25_can_lehmann_fsm__2911_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net966 sg13g2_dlygate4sd3_1
XFILLER_6_216 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_hold989 heichips25_can_lehmann_fsm/_0094_ VPWR VGND heichips25_can_lehmann_fsm/net988
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold978 heichips25_can_lehmann_fsm__2883_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net977 sg13g2_dlygate4sd3_1
Xheichips25_sap3__3750_ VPWR heichips25_sap3/_1262_ heichips25_sap3/net293 VGND sg13g2_inv_1
Xheichips25_sap3__3681_ heichips25_sap3/_0143_ heichips25_sap3/_1129_ heichips25_sap3/_1222_
+ heichips25_sap3/net111 heichips25_sap3/_1422_ VPWR VGND sg13g2_a22oi_1
XFILLER_40_98 VPWR VGND sg13g2_fill_2
XFILLER_3_956 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2701_ heichips25_sap3/net274 heichips25_sap3__3922_/Q heichips25_sap3/_0347_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__2632_ VGND VPWR heichips25_sap3/_1503_ heichips25_sap3/_1568_ heichips25_sap3/_0299_
+ heichips25_sap3/_0295_ sg13g2_a21oi_1
Xheichips25_sap3__2563_ heichips25_sap3/_0238_ heichips25_sap3/net73 heichips25_sap3__4006_/Q
+ heichips25_sap3/net81 heichips25_sap3__3974_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2494_ heichips25_sap3/_1902_ heichips25_sap3/_1903_ heichips25_sap3/_1905_
+ heichips25_sap3/_1906_ heichips25_sap3/_1907_ VPWR VGND sg13g2_and4_1
XFILLER_18_334 VPWR VGND sg13g2_decap_8
XFILLER_19_846 VPWR VGND sg13g2_fill_2
XFILLER_46_654 VPWR VGND sg13g2_decap_8
XFILLER_18_356 VPWR VGND sg13g2_fill_2
XFILLER_34_849 VPWR VGND sg13g2_decap_4
XFILLER_45_197 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3115_ heichips25_sap3/_1719_ heichips25_sap3/_0698_ heichips25_sap3/_0725_
+ heichips25_sap3/_0727_ heichips25_sap3/_0728_ VPWR VGND sg13g2_or4_1
Xheichips25_sap3__3046_ heichips25_sap3/_0658_ VPWR heichips25_sap3/_0659_ VGND heichips25_sap3/_0640_
+ heichips25_sap3/_0653_ sg13g2_o21ai_1
Xheichips25_sap3__3948_ heichips25_sap3/net433 VGND VPWR heichips25_sap3/_0089_ heichips25_sap3__3948_/Q
+ heichips25_sap3__3996_/CLK sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1982_ heichips25_can_lehmann_fsm/_0334_ heichips25_can_lehmann_fsm__2783_/Q
+ heichips25_can_lehmann_fsm/_0340_ VPWR VGND sg13g2_nor2b_1
XFILLER_49_492 VPWR VGND sg13g2_fill_2
Xinput3 ui_in[0] net3 VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm__2603_ VGND VPWR heichips25_can_lehmann_fsm/_0897_ heichips25_can_lehmann_fsm/net422
+ heichips25_can_lehmann_fsm/_0201_ heichips25_can_lehmann_fsm/_0767_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2534_ heichips25_can_lehmann_fsm/net476 VPWR heichips25_can_lehmann_fsm/_0733_
+ VGND heichips25_can_lehmann_fsm__2942_/Q heichips25_can_lehmann_fsm/net395 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2465_ VGND VPWR heichips25_can_lehmann_fsm/_0931_ heichips25_can_lehmann_fsm/net386
+ heichips25_can_lehmann_fsm/_0132_ heichips25_can_lehmann_fsm/_0698_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2396_ heichips25_can_lehmann_fsm/net470 VPWR heichips25_can_lehmann_fsm/_0664_
+ VGND heichips25_can_lehmann_fsm__2873_/Q heichips25_can_lehmann_fsm/net390 sg13g2_o21ai_1
XFILLER_10_57 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__3017_ net746 VGND VPWR heichips25_can_lehmann_fsm/net999
+ heichips25_can_lehmann_fsm__3017_/Q clknet_leaf_20_clk sg13g2_dfrbpq_1
XFILLER_0_915 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2790__627 VPWR VGND net626 sg13g2_tiehi
XFILLER_27_131 VPWR VGND sg13g2_decap_8
XFILLER_15_304 VPWR VGND sg13g2_fill_1
XFILLER_16_827 VPWR VGND sg13g2_fill_2
XFILLER_16_849 VPWR VGND sg13g2_fill_2
XFILLER_28_687 VPWR VGND sg13g2_fill_2
XFILLER_24_871 VPWR VGND sg13g2_decap_4
XFILLER_42_189 VPWR VGND sg13g2_decap_8
XFILLER_23_370 VPWR VGND sg13g2_decap_8
XFILLER_11_543 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3802_ heichips25_sap3/net340 heichips25_sap3/net925 heichips25_sap3/_1310_
+ heichips25_sap3/_0176_ VPWR VGND sg13g2_a21o_1
Xheichips25_sap3__1994_ VPWR heichips25_sap3/_1420_ heichips25_sap3__3938_/Q VGND
+ sg13g2_inv_1
XFILLER_3_731 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3733_ heichips25_sap3/_1249_ VPWR heichips25_sap3/_1250_ VGND heichips25_sap3__4029_/Q
+ heichips25_sap3/net1011 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2836__535 VPWR VGND net534 sg13g2_tiehi
XFILLER_3_764 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3664_ heichips25_sap3/net146 VPWR heichips25_sap3/_1209_ VGND uio_oe_sap3\[4\]
+ heichips25_sap3/_0732_ sg13g2_o21ai_1
Xheichips25_sap3__3595_ uio_oe_sap3\[7\] net47 heichips25_sap3/_1144_ heichips25_sap3/_1169_
+ VPWR VGND sg13g2_mux2_1
Xheichips25_sap3__2615_ heichips25_sap3/_1592_ VPWR heichips25_sap3__4070_/A VGND
+ heichips25_sap3/_1471_ heichips25_sap3/_0285_ sg13g2_o21ai_1
Xheichips25_sap3__2546_ heichips25_sap3/net215 heichips25_sap3/_0221_ heichips25_sap3/_0222_
+ VPWR VGND sg13g2_nor2_1
XFILLER_19_610 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2477_ VGND VPWR heichips25_sap3/net265 heichips25_sap3/_1879_ heichips25_sap3/_1890_
+ heichips25_sap3/net212 sg13g2_a21oi_1
XFILLER_18_175 VPWR VGND sg13g2_decap_8
XFILLER_15_871 VPWR VGND sg13g2_fill_2
XFILLER_21_318 VPWR VGND sg13g2_fill_2
XFILLER_30_830 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3029_ heichips25_sap3/_1521_ heichips25_sap3/_1527_ heichips25_sap3/_1504_
+ heichips25_sap3/_0642_ VPWR VGND heichips25_sap3/_1565_ sg13g2_nand4_1
XFILLER_30_852 VPWR VGND sg13g2_decap_4
XFILLER_30_863 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2250_ heichips25_can_lehmann_fsm/_0570_ heichips25_can_lehmann_fsm/net1173
+ heichips25_can_lehmann_fsm/_1043_ VPWR VGND sg13g2_nand2b_1
Xheichips25_can_lehmann_fsm__2181_ heichips25_can_lehmann_fsm/_0516_ heichips25_can_lehmann_fsm/net164
+ heichips25_can_lehmann_fsm/_0515_ VPWR VGND sg13g2_nand2_1
Xheichips25_can_lehmann_fsm__1965_ VPWR VGND heichips25_can_lehmann_fsm/net192 heichips25_can_lehmann_fsm/_0325_
+ heichips25_can_lehmann_fsm/_0324_ heichips25_can_lehmann_fsm/_0322_ heichips25_can_lehmann_fsm/_0005_
+ heichips25_can_lehmann_fsm/_0323_ sg13g2_a221oi_1
XFILLER_38_996 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1896_ heichips25_can_lehmann_fsm/_1209_ heichips25_can_lehmann_fsm/net307
+ heichips25_can_lehmann_fsm__2953_/Q heichips25_can_lehmann_fsm/net311 heichips25_can_lehmann_fsm__3025_/Q
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3_hold1113 heichips25_sap3__4056_/Q VPWR VGND heichips25_sap3/net1112
+ sg13g2_dlygate4sd3_1
XFILLER_13_808 VPWR VGND sg13g2_fill_1
Xheichips25_sap3_hold1146 heichips25_sap3__4049_/Q VPWR VGND heichips25_sap3/net1145
+ sg13g2_dlygate4sd3_1
Xheichips25_sap3_hold1179 heichips25_sap3__4041_/Q VPWR VGND heichips25_sap3/net1178
+ sg13g2_dlygate4sd3_1
XFILLER_33_690 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2517_ VGND VPWR heichips25_can_lehmann_fsm/_0918_ heichips25_can_lehmann_fsm/net378
+ heichips25_can_lehmann_fsm/_0158_ heichips25_can_lehmann_fsm/_0724_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2448_ heichips25_can_lehmann_fsm/net468 VPWR heichips25_can_lehmann_fsm/_0690_
+ VGND heichips25_can_lehmann_fsm__2898_/Q heichips25_can_lehmann_fsm/net359 sg13g2_o21ai_1
XFILLER_4_506 VPWR VGND sg13g2_fill_1
XFILLER_20_395 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2379_ VGND VPWR heichips25_can_lehmann_fsm/_0957_ heichips25_can_lehmann_fsm/net423
+ heichips25_can_lehmann_fsm/_0089_ heichips25_can_lehmann_fsm/_0655_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm_fanout472 heichips25_can_lehmann_fsm/net474 heichips25_can_lehmann_fsm/net472
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout483 heichips25_can_lehmann_fsm/net484 heichips25_can_lehmann_fsm/net483
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout494 heichips25_can_lehmann_fsm/net496 heichips25_can_lehmann_fsm/net494
+ VPWR VGND sg13g2_buf_1
XFILLER_43_1014 VPWR VGND sg13g2_fill_2
XFILLER_0_745 VPWR VGND sg13g2_fill_1
XFILLER_43_1025 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2400_ heichips25_sap3/_1819_ heichips25_sap3/net73 heichips25_sap3__4009_/Q
+ heichips25_sap3/net81 heichips25_sap3__3977_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_47_215 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3380_ heichips25_sap3/_0988_ heichips25_sap3/net132 heichips25_sap3__3992_/Q
+ heichips25_sap3/net135 heichips25_sap3__3968_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2331_ VPWR VGND heichips25_sap3/_1751_ heichips25_sap3/_1654_ heichips25_sap3/_1747_
+ heichips25_sap3/_1420_ heichips25_sap3/_1752_ heichips25_sap3/net90 sg13g2_a221oi_1
XFILLER_46_53 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2262_ heichips25_sap3/_1544_ heichips25_sap3/_1553_ heichips25_sap3/net229
+ heichips25_sap3/_1683_ VPWR VGND heichips25_sap3/_1681_ sg13g2_nand4_1
XFILLER_44_944 VPWR VGND sg13g2_decap_4
XFILLER_43_421 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__4001_ heichips25_sap3/net440 VGND VPWR heichips25_sap3/_0142_ heichips25_sap3__4001_/Q
+ heichips25_sap3__4018_/CLK sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2946__552 VPWR VGND net551 sg13g2_tiehi
XFILLER_44_988 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2193_ heichips25_sap3__3929_/Q heichips25_sap3/net259 heichips25_sap3/_1614_
+ VPWR VGND sg13g2_nor2b_1
XFILLER_15_178 VPWR VGND sg13g2_fill_1
XFILLER_31_638 VPWR VGND sg13g2_fill_2
XFILLER_7_333 VPWR VGND sg13g2_fill_2
XFILLER_7_322 VPWR VGND sg13g2_decap_8
XFILLER_8_845 VPWR VGND sg13g2_fill_1
XFILLER_7_69 VPWR VGND sg13g2_fill_1
XFILLER_7_58 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__1977_ VPWR heichips25_sap3/_1403_ heichips25_sap3__3983_/Q VGND
+ sg13g2_inv_1
Xheichips25_sap3__3716_ heichips25_sap3/_0159_ heichips25_sap3/_1129_ heichips25_sap3/_1241_
+ heichips25_sap3/net114 heichips25_sap3/_1421_ VPWR VGND sg13g2_a22oi_1
XFILLER_39_705 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3647_ heichips25_sap3/_1195_ VPWR heichips25_sap3/_1196_ VGND heichips25_sap3/_0777_
+ heichips25_sap3/_0870_ sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2888__720 VPWR VGND net719 sg13g2_tiehi
Xheichips25_sap3__3578_ uio_oe_sap3\[3\] heichips25_sap3/net95 heichips25_sap3/_1156_
+ VPWR VGND sg13g2_nor2_1
XFILLER_38_248 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2529_ heichips25_sap3/_0204_ heichips25_sap3/_0205_ heichips25_sap3/_0206_
+ VPWR VGND sg13g2_and2_1
Xheichips25_can_lehmann_fsm__1750_ VGND VPWR heichips25_can_lehmann_fsm/_1070_ heichips25_can_lehmann_fsm/_1069_
+ heichips25_can_lehmann_fsm/_1068_ sg13g2_or2_1
Xheichips25_can_lehmann_fsm__1681_ heichips25_can_lehmann_fsm/_1005_ heichips25_can_lehmann_fsm/net296
+ heichips25_can_lehmann_fsm__2897_/Q heichips25_can_lehmann_fsm/net317 heichips25_can_lehmann_fsm__2993_/Q
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2925__636 VPWR VGND net635 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2302_ heichips25_can_lehmann_fsm/_1052_ heichips25_can_lehmann_fsm/_0611_
+ heichips25_can_lehmann_fsm/_0612_ VPWR VGND sg13g2_nor2b_1
Xheichips25_can_lehmann_fsm__2233_ VGND VPWR heichips25_can_lehmann_fsm/net161 heichips25_can_lehmann_fsm/_0555_
+ heichips25_can_lehmann_fsm/_0042_ heichips25_can_lehmann_fsm/_0556_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2164_ heichips25_can_lehmann_fsm/_0502_ heichips25_can_lehmann_fsm/net1233
+ heichips25_can_lehmann_fsm/net1226 VPWR VGND sg13g2_xnor2_1
Xheichips25_can_lehmann_fsm__2095_ VGND VPWR heichips25_can_lehmann_fsm/_0434_ heichips25_can_lehmann_fsm/_0435_
+ heichips25_can_lehmann_fsm/_0024_ heichips25_can_lehmann_fsm/_0436_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2997_ net617 VGND VPWR heichips25_can_lehmann_fsm/_0222_
+ heichips25_can_lehmann_fsm__2997_/Q clknet_leaf_0_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1948_ heichips25_can_lehmann_fsm/_0311_ heichips25_can_lehmann_fsm/net186
+ heichips25_can_lehmann_fsm/_0310_ heichips25_can_lehmann_fsm/net199 heichips25_can_lehmann_fsm/net1262
+ VPWR VGND sg13g2_a22oi_1
XFILLER_38_793 VPWR VGND sg13g2_fill_1
XFILLER_26_922 VPWR VGND sg13g2_decap_8
XFILLER_26_966 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1879_ heichips25_can_lehmann_fsm/_1190_ heichips25_can_lehmann_fsm/_1191_
+ heichips25_can_lehmann_fsm/_1189_ heichips25_can_lehmann_fsm/_1193_ VPWR VGND heichips25_can_lehmann_fsm/_1192_
+ sg13g2_nand4_1
XFILLER_12_137 VPWR VGND sg13g2_decap_8
XFILLER_5_804 VPWR VGND sg13g2_fill_2
XFILLER_20_181 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2880_ heichips25_sap3/_0521_ heichips25_sap3/_0445_ heichips25_sap3/_0356_
+ heichips25_sap3/_0406_ heichips25_sap3/net154 VPWR VGND sg13g2_a22oi_1
XFILLER_4_358 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3501_ uio_out_sap3\[1\] heichips25_sap3/net131 heichips25_sap3/_1097_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__3432_ heichips25_sap3/_1038_ heichips25_sap3/net54 heichips25_sap3/_0873_
+ VPWR VGND sg13g2_xnor2_1
Xheichips25_sap3__3363_ VGND VPWR heichips25_sap3/_0820_ heichips25_sap3/_0934_ heichips25_sap3/_0972_
+ heichips25_sap3/net63 sg13g2_a21oi_1
XFILLER_35_229 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2314_ heichips25_sap3/_1680_ heichips25_sap3/_1693_ heichips25_sap3/_1712_
+ heichips25_sap3/_1732_ heichips25_sap3/_1735_ VPWR VGND sg13g2_nor4_1
Xheichips25_sap3__3294_ heichips25_sap3/_0906_ heichips25_sap3/_1922_ heichips25_sap3/_0884_
+ VPWR VGND sg13g2_nand2_1
XFILLER_28_292 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2245_ heichips25_sap3/_1537_ heichips25_sap3/_1551_ heichips25_sap3/_1459_
+ heichips25_sap3/_1666_ VPWR VGND sg13g2_nand3_1
XFILLER_43_295 VPWR VGND sg13g2_fill_1
XFILLER_43_262 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2176_ heichips25_sap3/_1478_ heichips25_sap3/_1567_ heichips25_sap3/_1597_
+ VPWR VGND sg13g2_nor2_1
XFILLER_31_468 VPWR VGND sg13g2_fill_2
XFILLER_8_642 VPWR VGND sg13g2_fill_2
XFILLER_4_870 VPWR VGND sg13g2_decap_8
XFILLER_39_535 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2920_ net655 VGND VPWR heichips25_can_lehmann_fsm/net982
+ heichips25_can_lehmann_fsm__2920_/Q clknet_leaf_19_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2851_ net793 VGND VPWR heichips25_can_lehmann_fsm/_0076_
+ heichips25_can_lehmann_fsm__2851_/Q clknet_leaf_8_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1802_ heichips25_can_lehmann_fsm/net337 VPWR heichips25_can_lehmann_fsm/_1118_
+ VGND heichips25_can_lehmann_fsm__2972_/Q heichips25_can_lehmann_fsm/net338 sg13g2_o21ai_1
XFILLER_26_218 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2782_ net642 VGND VPWR heichips25_can_lehmann_fsm/net1258
+ heichips25_can_lehmann_fsm__2782_/Q clknet_leaf_5_clk sg13g2_dfrbpq_1
Xheichips25_sap3_clk_div_param_inst_clock_root heichips25_sap3/clk_div_out heichips25_sap3_clk_div_param_inst__2_/Q
+ VPWR VGND sg13g2_buf_16
Xheichips25_can_lehmann_fsm__1733_ heichips25_can_lehmann_fsm/_1054_ heichips25_can_lehmann_fsm/_1053_
+ heichips25_can_lehmann_fsm/_1051_ VPWR VGND sg13g2_nand2b_1
XFILLER_22_435 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1664_ VPWR heichips25_can_lehmann_fsm/_0988_ net6 VGND
+ sg13g2_inv_1
Xheichips25_can_lehmann_fsm__1595_ VPWR heichips25_can_lehmann_fsm/_0919_ heichips25_can_lehmann_fsm/net992
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__2216_ VGND VPWR heichips25_can_lehmann_fsm/net162 heichips25_can_lehmann_fsm/_0542_
+ heichips25_can_lehmann_fsm/_0038_ heichips25_can_lehmann_fsm/_0543_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2147_ heichips25_can_lehmann_fsm/_0485_ VPWR heichips25_can_lehmann_fsm/_0486_
+ VGND heichips25_can_lehmann_fsm/_0884_ heichips25_can_lehmann_fsm/_0991_ sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2078_ VGND VPWR heichips25_can_lehmann_fsm/_0417_ heichips25_can_lehmann_fsm/_0421_
+ heichips25_can_lehmann_fsm/_0021_ heichips25_can_lehmann_fsm/_0422_ sg13g2_a21oi_1
XFILLER_27_44 VPWR VGND sg13g2_decap_8
XFILLER_38_590 VPWR VGND sg13g2_fill_2
XFILLER_41_700 VPWR VGND sg13g2_decap_8
Xheichips25_sap3_fanout140 heichips25_sap3/net141 heichips25_sap3/net140 VPWR VGND
+ sg13g2_buf_1
XFILLER_27_88 VPWR VGND sg13g2_fill_2
XFILLER_43_32 VPWR VGND sg13g2_decap_8
XFILLER_41_711 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2030_ heichips25_sap3/_1448_ heichips25_sap3/_1450_ heichips25_sap3/_1451_
+ VPWR VGND sg13g2_nor2_1
XFILLER_13_424 VPWR VGND sg13g2_fill_2
Xheichips25_sap3_fanout151 heichips25_sap3/_0751_ heichips25_sap3/net151 VPWR VGND
+ sg13g2_buf_1
XFILLER_13_446 VPWR VGND sg13g2_decap_8
XFILLER_13_457 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm_hold1230 heichips25_can_lehmann_fsm__3044_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1229 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1241 heichips25_can_lehmann_fsm__2787_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1240 sg13g2_dlygate4sd3_1
XFILLER_43_76 VPWR VGND sg13g2_fill_2
XFILLER_41_788 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm_hold1263 heichips25_can_lehmann_fsm__2793_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1262 sg13g2_dlygate4sd3_1
XFILLER_40_276 VPWR VGND sg13g2_fill_2
XFILLER_40_265 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm_hold1252 heichips25_can_lehmann_fsm__2785_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1251 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1274 heichips25_can_lehmann_fsm__2776_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1273 sg13g2_dlygate4sd3_1
Xclkbuf_leaf_20_clk clknet_2_2__leaf_clk clknet_leaf_20_clk VPWR VGND sg13g2_buf_8
Xheichips25_sap3__3981_ heichips25_sap3/net434 VGND VPWR heichips25_sap3/_0122_ heichips25_sap3__3981_/Q
+ heichips25_sap3__4012_/CLK sg13g2_dfrbpq_1
Xheichips25_sap3__2932_ VPWR VGND heichips25_sap3/_1384_ heichips25_sap3/_0570_ heichips25_sap3/_0442_
+ heichips25_sap3/_0343_ heichips25_sap3/_0571_ heichips25_sap3/_0399_ sg13g2_a221oi_1
Xheichips25_sap3__2863_ heichips25_sap3/_0505_ heichips25_sap3/_0504_ heichips25_sap3/_0501_
+ VPWR VGND sg13g2_nand2b_1
Xheichips25_sap3__2794_ heichips25_sap3/_1897_ heichips25_sap3/_0438_ heichips25_sap3/_1885_
+ heichips25_sap3/_0439_ VPWR VGND sg13g2_nand3_1
XFILLER_4_37 VPWR VGND sg13g2_decap_4
XFILLER_4_26 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3415_ VGND VPWR heichips25_sap3/net123 heichips25_sap3/_1021_ heichips25_sap3/_1022_
+ heichips25_sap3/_0863_ sg13g2_a21oi_1
Xheichips25_sap3__3346_ VGND VPWR heichips25_sap3/net45 heichips25_sap3/_0884_ heichips25_sap3/_0956_
+ heichips25_sap3/_0955_ sg13g2_a21oi_1
XFILLER_16_240 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3277_ heichips25_sap3/_0861_ heichips25_sap3/_0876_ heichips25_sap3/_0747_
+ heichips25_sap3/_0890_ VPWR VGND heichips25_sap3/_0887_ sg13g2_nand4_1
Xheichips25_sap3__2228_ heichips25_sap3/_1450_ heichips25_sap3/_1616_ heichips25_sap3/_1649_
+ VPWR VGND sg13g2_nor2_1
XFILLER_32_755 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2159_ heichips25_sap3/_1580_ heichips25_sap3/_1551_ heichips25_sap3/_1566_
+ heichips25_sap3/_1546_ heichips25_sap3/_1463_ VPWR VGND sg13g2_a22oi_1
XFILLER_20_939 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_11_clk clknet_2_3__leaf_clk clknet_leaf_11_clk VPWR VGND sg13g2_buf_8
XFILLER_9_995 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__3050_ net541 VGND VPWR heichips25_can_lehmann_fsm/net1118
+ heichips25_can_lehmann_fsm__3050_/Q clknet_leaf_12_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2001_ VGND VPWR heichips25_can_lehmann_fsm/net180 heichips25_can_lehmann_fsm/_0355_
+ heichips25_can_lehmann_fsm/_0010_ heichips25_can_lehmann_fsm/_0356_ sg13g2_a21oi_1
XFILLER_39_321 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2903_ net689 VGND VPWR heichips25_can_lehmann_fsm/_0128_
+ heichips25_can_lehmann_fsm__2903_/Q clknet_leaf_6_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2834_ net538 VGND VPWR heichips25_can_lehmann_fsm/_0059_
+ heichips25_can_lehmann_fsm__2834_/Q clknet_leaf_5_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2765_ VGND VPWR heichips25_can_lehmann_fsm/_0853_ heichips25_can_lehmann_fsm/net375
+ heichips25_can_lehmann_fsm/_0282_ heichips25_can_lehmann_fsm/_0848_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__1716_ VGND VPWR heichips25_can_lehmann_fsm/net1277 heichips25_can_lehmann_fsm/_1016_
+ heichips25_can_lehmann_fsm/_1039_ heichips25_can_lehmann_fsm/_1029_ sg13g2_a21oi_1
XFILLER_23_733 VPWR VGND sg13g2_fill_1
Xfanout47 net47 uio_out_sap3\[7\] VPWR VGND sg13g2_buf_4
Xheichips25_can_lehmann_fsm__2696_ heichips25_can_lehmann_fsm/net475 VPWR heichips25_can_lehmann_fsm/_0814_
+ VGND heichips25_can_lehmann_fsm__3023_/Q heichips25_can_lehmann_fsm/net406 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__1647_ VPWR heichips25_can_lehmann_fsm/_0971_ heichips25_can_lehmann_fsm/net1093
+ VGND sg13g2_inv_1
XFILLER_10_416 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1578_ VPWR heichips25_can_lehmann_fsm/_0902_ heichips25_can_lehmann_fsm/net874
+ VGND sg13g2_inv_1
XFILLER_13_35 VPWR VGND sg13g2_fill_2
XFILLER_13_46 VPWR VGND sg13g2_decap_8
XFILLER_1_125 VPWR VGND sg13g2_decap_8
XFILLER_38_65 VPWR VGND sg13g2_fill_1
XFILLER_18_538 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3200_ heichips25_sap3/_0813_ heichips25_sap3/net138 heichips25_sap3__3982_/Q
+ heichips25_sap3/net140 heichips25_sap3__3990_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_45_368 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3131_ heichips25_sap3/_0656_ VPWR heichips25_sap3/_0744_ VGND heichips25_sap3/_0435_
+ heichips25_sap3/_0743_ sg13g2_o21ai_1
XFILLER_14_711 VPWR VGND sg13g2_fill_2
XFILLER_14_722 VPWR VGND sg13g2_decap_4
XFILLER_41_541 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3062_ heichips25_sap3/_0673_ heichips25_sap3/_0674_ heichips25_sap3/_0672_
+ heichips25_sap3/_0675_ VPWR VGND sg13g2_nand3_1
XFILLER_41_574 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2013_ heichips25_sap3/net258 heichips25_sap3/net260 heichips25_sap3/_1434_
+ VPWR VGND sg13g2_nor2_1
XFILLER_9_214 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm_hold1071 heichips25_can_lehmann_fsm__2918_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1070 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1082 heichips25_can_lehmann_fsm__2870_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1081 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1093 heichips25_can_lehmann_fsm__2926_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1092 sg13g2_dlygate4sd3_1
XFILLER_10_950 VPWR VGND sg13g2_fill_1
Xclkload17 clknet_leaf_12_clk clkload17/X VPWR VGND sg13g2_buf_8
Xheichips25_sap3__3964_ heichips25_sap3/net434 VGND VPWR heichips25_sap3/_0105_ heichips25_sap3__3964_/Q
+ heichips25_sap3__3996_/CLK sg13g2_dfrbpq_1
Xclkload28 VPWR clkload28/Y clkload28/A VGND sg13g2_inv_1
Xheichips25_sap3__2915_ heichips25_sap3/_0555_ heichips25_sap3/_0552_ heichips25_sap3/_0554_
+ VPWR VGND sg13g2_xnor2_1
Xheichips25_sap3__3895_ heichips25_sap3/net448 VGND VPWR heichips25_sap3/_0036_ heichips25_sap3__3895_/Q
+ net819 sg13g2_dfrbpq_1
XFILLER_5_486 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2846_ heichips25_sap3/_0375_ heichips25_sap3/_0374_ heichips25_sap3/_0489_
+ VPWR VGND sg13g2_xor2_1
Xheichips25_can_lehmann_fsm__3017__747 VPWR VGND net746 sg13g2_tiehi
Xheichips25_sap3__2777_ VGND VPWR heichips25_sap3/_1880_ heichips25_sap3/_0420_ heichips25_sap3/_0423_
+ heichips25_sap3/_0422_ sg13g2_a21oi_1
Xclkbuf_leaf_0_clk clknet_2_0__leaf_clk clknet_leaf_0_clk VPWR VGND sg13g2_buf_8
XFILLER_49_696 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3329_ heichips25_sap3/_0939_ heichips25_sap3/net133 heichips25_sap3__3990_/Q
+ heichips25_sap3/net137 heichips25_sap3__3966_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2550_ heichips25_can_lehmann_fsm/net473 VPWR heichips25_can_lehmann_fsm/_0741_
+ VGND heichips25_can_lehmann_fsm__2950_/Q heichips25_can_lehmann_fsm/net402 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2481_ VGND VPWR heichips25_can_lehmann_fsm/_0927_ heichips25_can_lehmann_fsm/net370
+ heichips25_can_lehmann_fsm/_0140_ heichips25_can_lehmann_fsm/_0706_ sg13g2_a21oi_1
XFILLER_9_770 VPWR VGND sg13g2_fill_1
Xclkbuf_5_31__f_heichips25_sap3\_sap_3_inst.alu_inst.clk clkload29/A clknet_4_15_0_heichips25_sap3\/sap_3_inst.alu_inst.clk
+ VPWR VGND sg13g2_buf_16
Xheichips25_can_lehmann_fsm__3033_ net581 VGND VPWR heichips25_can_lehmann_fsm/net994
+ heichips25_can_lehmann_fsm__3033_/Q clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_5_91 VPWR VGND sg13g2_decap_4
XFILLER_8_1028 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__3033__582 VPWR VGND net581 sg13g2_tiehi
XFILLER_27_302 VPWR VGND sg13g2_decap_8
XFILLER_39_195 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2817_ net572 VGND VPWR heichips25_can_lehmann_fsm/net1206
+ heichips25_can_lehmann_fsm__2817_/Q clknet_leaf_7_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2748_ heichips25_can_lehmann_fsm/net491 VPWR heichips25_can_lehmann_fsm/_0840_
+ VGND heichips25_can_lehmann_fsm/net1127 heichips25_can_lehmann_fsm/net380 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm_hold913 heichips25_can_lehmann_fsm__2866_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net912 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold924 heichips25_can_lehmann_fsm__3012_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net923 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__2679_ VGND VPWR heichips25_can_lehmann_fsm/_0876_ heichips25_can_lehmann_fsm/net395
+ heichips25_can_lehmann_fsm/_0239_ heichips25_can_lehmann_fsm/_0805_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm_hold935 heichips25_can_lehmann_fsm__2947_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net934 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold902 heichips25_can_lehmann_fsm/_0132_ VPWR VGND heichips25_can_lehmann_fsm/net901
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold957 heichips25_can_lehmann_fsm/_0116_ VPWR VGND heichips25_can_lehmann_fsm/net956
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold946 heichips25_can_lehmann_fsm/_0265_ VPWR VGND heichips25_can_lehmann_fsm/net945
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold968 heichips25_can_lehmann_fsm/_0136_ VPWR VGND heichips25_can_lehmann_fsm/net967
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold979 heichips25_can_lehmann_fsm__2985_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net978 sg13g2_dlygate4sd3_1
XFILLER_3_913 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3680_ VGND VPWR heichips25_sap3/_0888_ heichips25_sap3/_1220_ heichips25_sap3/_1222_
+ heichips25_sap3/_1221_ sg13g2_a21oi_1
XFILLER_3_946 VPWR VGND sg13g2_fill_1
XFILLER_3_924 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2700_ heichips25_sap3/_0346_ heichips25_sap3/_0339_ heichips25_sap3/_0345_
+ VPWR VGND sg13g2_nand2_1
XFILLER_2_423 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2631_ heichips25_sap3/net244 heichips25_sap3/_1551_ heichips25_sap3/_1459_
+ heichips25_sap3/_0298_ VPWR VGND sg13g2_nand3_1
XFILLER_49_53 VPWR VGND sg13g2_decap_8
XFILLER_49_75 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2562_ VPWR VGND heichips25_sap3__3982_/Q heichips25_sap3/net79 heichips25_sap3/net71
+ heichips25_sap3__3966_/Q heichips25_sap3/_0237_ heichips25_sap3/net83 sg13g2_a221oi_1
Xheichips25_sap3__2493_ heichips25_sap3/_1906_ heichips25_sap3/net82 heichips25_sap3__3964_/Q
+ heichips25_sap3/net83 heichips25_sap3__3956_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_18_313 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2847__802 VPWR VGND net801 sg13g2_tiehi
XFILLER_34_839 VPWR VGND sg13g2_decap_4
XFILLER_33_327 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3114_ heichips25_sap3/_0726_ VPWR heichips25_sap3/_0727_ VGND heichips25_sap3/_1527_
+ heichips25_sap3/_1871_ sg13g2_o21ai_1
Xheichips25_sap3__3045_ VGND VPWR heichips25_sap3/net220 heichips25_sap3/_0657_ heichips25_sap3/_0658_
+ heichips25_sap3/net248 sg13g2_a21oi_1
XFILLER_14_563 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3947_ heichips25_sap3/net439 VGND VPWR heichips25_sap3/_0088_ heichips25_sap3__3947_/Q
+ heichips25_sap3__4015_/CLK sg13g2_dfrbpq_1
XFILLER_5_294 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2829_ heichips25_sap3/_0472_ VPWR heichips25_sap3/_0473_ VGND heichips25_sap3/net64
+ heichips25_sap3/_0471_ sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__1981_ heichips25_can_lehmann_fsm__2783_/Q heichips25_can_lehmann_fsm/_0334_
+ heichips25_can_lehmann_fsm/_0339_ VPWR VGND sg13g2_nor2b_1
XFILLER_49_471 VPWR VGND sg13g2_fill_2
Xinput4 ui_in[1] net4 VPWR VGND sg13g2_buf_1
Xclkbuf_2_1__f_clk clknet_2_1__leaf_clk clknet_0_clk VPWR VGND sg13g2_buf_16
XFILLER_36_176 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2602_ heichips25_can_lehmann_fsm/net493 VPWR heichips25_can_lehmann_fsm/_0767_
+ VGND heichips25_can_lehmann_fsm__2976_/Q heichips25_can_lehmann_fsm/net422 sg13g2_o21ai_1
XFILLER_17_390 VPWR VGND sg13g2_decap_8
XFILLER_33_850 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2533_ VGND VPWR heichips25_can_lehmann_fsm/_0914_ heichips25_can_lehmann_fsm/net368
+ heichips25_can_lehmann_fsm/_0166_ heichips25_can_lehmann_fsm/_0732_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2898__700 VPWR VGND net699 sg13g2_tiehi
XFILLER_32_393 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2464_ heichips25_can_lehmann_fsm/net499 VPWR heichips25_can_lehmann_fsm/_0698_
+ VGND heichips25_can_lehmann_fsm__2906_/Q heichips25_can_lehmann_fsm/net386 sg13g2_o21ai_1
XFILLER_20_555 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2395_ VGND VPWR heichips25_can_lehmann_fsm/_0953_ heichips25_can_lehmann_fsm/net390
+ heichips25_can_lehmann_fsm/_0097_ heichips25_can_lehmann_fsm/_0663_ sg13g2_a21oi_1
XFILLER_3_209 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__3016_ net754 VGND VPWR heichips25_can_lehmann_fsm/net854
+ heichips25_can_lehmann_fsm__3016_/Q clknet_leaf_19_clk sg13g2_dfrbpq_1
XFILLER_28_666 VPWR VGND sg13g2_fill_1
XFILLER_42_102 VPWR VGND sg13g2_decap_4
XFILLER_24_861 VPWR VGND sg13g2_fill_1
XFILLER_11_533 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3801_ VPWR VGND heichips25_sap3/_1309_ heichips25_sap3/net339 heichips25_sap3/_1303_
+ heichips25_sap3/_1368_ heichips25_sap3/_1310_ heichips25_sap3/net290 sg13g2_a221oi_1
Xheichips25_sap3__3732_ VGND VPWR heichips25_sap3__4029_/Q heichips25_sap3/_1426_
+ heichips25_sap3/_1249_ heichips25_sap3__4030_/Q sg13g2_a21oi_1
Xheichips25_sap3__1993_ VPWR heichips25_sap3/_1419_ heichips25_sap3__3945_/Q VGND
+ sg13g2_inv_1
XFILLER_2_253 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3663_ heichips25_sap3/_0139_ heichips25_sap3/_1106_ heichips25_sap3/_1208_
+ heichips25_sap3/net112 heichips25_sap3/_1370_ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3594_ heichips25_sap3/_0110_ heichips25_sap3/_1124_ heichips25_sap3/_1168_
+ heichips25_sap3/net101 heichips25_sap3/_1417_ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2614_ heichips25_sap3/_0280_ heichips25_sap3/_0283_ heichips25_sap3/_0284_
+ heichips25_sap3/_0285_ VPWR VGND sg13g2_nor3_1
Xheichips25_sap3__2545_ heichips25_sap3/_0220_ VPWR heichips25_sap3/_0221_ VGND heichips25_sap3/_0214_
+ heichips25_sap3/_0217_ sg13g2_o21ai_1
XFILLER_47_964 VPWR VGND sg13g2_fill_2
XFILLER_46_430 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2476_ heichips25_sap3/_1619_ heichips25_sap3/_1714_ heichips25_sap3/_1889_
+ VPWR VGND sg13g2_nor2_1
XFILLER_18_143 VPWR VGND sg13g2_decap_8
XFILLER_20_1026 VPWR VGND sg13g2_fill_2
XFILLER_46_474 VPWR VGND sg13g2_fill_1
XFILLER_34_669 VPWR VGND sg13g2_fill_2
XFILLER_22_809 VPWR VGND sg13g2_fill_1
XFILLER_33_146 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3028_ heichips25_sap3/_1520_ heichips25_sap3/_1658_ heichips25_sap3/_0641_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_can_lehmann_fsm__2180_ heichips25_can_lehmann_fsm/_0515_ heichips25_can_lehmann_fsm/net1236
+ heichips25_can_lehmann_fsm/_1098_ VPWR VGND sg13g2_xnor2_1
Xheichips25_sap3_clk_div_param_inst__2_ heichips25_sap3/net450 VGND VPWR heichips25_sap3_clk_div_param_inst__2_/D
+ heichips25_sap3_clk_div_param_inst__2_/Q clknet_leaf_23_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1964_ heichips25_can_lehmann_fsm/net322 VPWR heichips25_can_lehmann_fsm/_0325_
+ VGND heichips25_can_lehmann_fsm/net1249 heichips25_can_lehmann_fsm/net178 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__1895_ heichips25_can_lehmann_fsm/_1208_ heichips25_can_lehmann_fsm/_1207_
+ heichips25_can_lehmann_fsm/net337 heichips25_can_lehmann_fsm/net333 heichips25_can_lehmann_fsm__3049_/Q
+ VPWR VGND sg13g2_a22oi_1
XFILLER_37_496 VPWR VGND sg13g2_fill_1
XFILLER_36_1000 VPWR VGND sg13g2_fill_1
Xheichips25_sap3_hold1125 heichips25_sap3__4054_/Q VPWR VGND heichips25_sap3/net1124
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__2516_ heichips25_can_lehmann_fsm/net485 VPWR heichips25_can_lehmann_fsm/_0724_
+ VGND heichips25_can_lehmann_fsm/net950 heichips25_can_lehmann_fsm/net378 sg13g2_o21ai_1
XFILLER_33_680 VPWR VGND sg13g2_fill_1
XFILLER_21_875 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2447_ VGND VPWR heichips25_can_lehmann_fsm/_0936_ heichips25_can_lehmann_fsm/net398
+ heichips25_can_lehmann_fsm/_0123_ heichips25_can_lehmann_fsm/_0689_ sg13g2_a21oi_1
XFILLER_21_897 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2378_ heichips25_can_lehmann_fsm/net495 VPWR heichips25_can_lehmann_fsm/_0655_
+ VGND heichips25_can_lehmann_fsm__2864_/Q heichips25_can_lehmann_fsm/net423 sg13g2_o21ai_1
XFILLER_21_79 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm_fanout473 heichips25_can_lehmann_fsm/net474 heichips25_can_lehmann_fsm/net473
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout484 heichips25_can_lehmann_fsm/net490 heichips25_can_lehmann_fsm/net484
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout495 heichips25_can_lehmann_fsm/net496 heichips25_can_lehmann_fsm/net495
+ VPWR VGND sg13g2_buf_1
Xheichips25_sap3__2330_ heichips25_sap3/_1738_ heichips25_sap3/_1748_ heichips25_sap3/_1749_
+ heichips25_sap3/_1750_ heichips25_sap3/_1751_ VPWR VGND sg13g2_and4_1
Xheichips25_sap3__2261_ VPWR heichips25_sap3/_1682_ heichips25_sap3/_1681_ VGND sg13g2_inv_1
XFILLER_28_485 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__4000_ heichips25_sap3/net440 VGND VPWR heichips25_sap3/_0141_ heichips25_sap3__4000_/Q
+ heichips25_sap3__4016_/CLK sg13g2_dfrbpq_1
Xheichips25_sap3__2192_ heichips25_sap3/net273 heichips25_sap3/net270 heichips25_sap3/net268
+ heichips25_sap3/_1613_ VPWR VGND sg13g2_nand3_1
XFILLER_31_606 VPWR VGND sg13g2_decap_4
XFILLER_30_127 VPWR VGND sg13g2_decap_4
XFILLER_7_356 VPWR VGND sg13g2_decap_8
XFILLER_8_879 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__1976_ VPWR heichips25_sap3/_1402_ heichips25_sap3__4007_/Q VGND
+ sg13g2_inv_1
Xheichips25_sap3__3715_ uio_oe_sap3\[7\] heichips25_sap3/net114 heichips25_sap3/_1131_
+ heichips25_sap3/_1241_ VPWR VGND sg13g2_nor3_1
Xheichips25_sap3__3646_ heichips25_sap3/net49 heichips25_sap3/_0889_ heichips25_sap3/_1195_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__3577_ heichips25_sap3/_0106_ heichips25_sap3/_0929_ heichips25_sap3/_1155_
+ heichips25_sap3/net100 heichips25_sap3/_1379_ VPWR VGND sg13g2_a22oi_1
XFILLER_19_430 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2528_ heichips25_sap3/_0205_ heichips25_sap3/net74 heichips25_sap3__4003_/Q
+ heichips25_sap3/net88 heichips25_sap3__3947_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2459_ heichips25_sap3/_1518_ heichips25_sap3/_1871_ heichips25_sap3/_1872_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_can_lehmann_fsm__1680_ heichips25_can_lehmann_fsm/net338 heichips25_can_lehmann_fsm/_0999_
+ heichips25_can_lehmann_fsm/_1004_ VPWR VGND sg13g2_nor2_1
XFILLER_34_433 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2301_ heichips25_can_lehmann_fsm/net1158 VPWR heichips25_can_lehmann_fsm/_0611_
+ VGND heichips25_can_lehmann_fsm__2830_/Q heichips25_can_lehmann_fsm/_1051_ sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2232_ heichips25_can_lehmann_fsm/net326 VPWR heichips25_can_lehmann_fsm/_0556_
+ VGND heichips25_can_lehmann_fsm/net1205 heichips25_can_lehmann_fsm/net161 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2163_ VPWR VGND heichips25_can_lehmann_fsm/_0501_ heichips25_can_lehmann_fsm/_1176_
+ heichips25_can_lehmann_fsm/_0500_ heichips25_can_lehmann_fsm/_0975_ heichips25_can_lehmann_fsm/_0027_
+ heichips25_can_lehmann_fsm/_0497_ sg13g2_a221oi_1
Xheichips25_can_lehmann_fsm__2094_ heichips25_can_lehmann_fsm/net322 VPWR heichips25_can_lehmann_fsm/_0436_
+ VGND heichips25_can_lehmann_fsm__2799_/Q heichips25_can_lehmann_fsm/net179 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2932__608 VPWR VGND net607 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2996_ net625 VGND VPWR heichips25_can_lehmann_fsm/_0221_
+ heichips25_can_lehmann_fsm__2996_/Q clknet_leaf_21_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1947_ heichips25_can_lehmann_fsm/_1061_ heichips25_can_lehmann_fsm/net1242
+ heichips25_can_lehmann_fsm/_0310_ VPWR VGND sg13g2_xor2_1
XFILLER_37_282 VPWR VGND sg13g2_fill_2
XFILLER_37_271 VPWR VGND sg13g2_decap_8
XFILLER_41_926 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1878_ VGND VPWR heichips25_can_lehmann_fsm__2892_/Q heichips25_can_lehmann_fsm/net297
+ heichips25_can_lehmann_fsm/_1192_ heichips25_can_lehmann_fsm/net302 sg13g2_a21oi_1
XFILLER_13_606 VPWR VGND sg13g2_fill_1
XFILLER_16_79 VPWR VGND sg13g2_fill_2
XFILLER_25_477 VPWR VGND sg13g2_decap_8
XFILLER_25_499 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3500_ heichips25_sap3/_1096_ heichips25_sap3/_0737_ heichips25_sap3/_1088_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__3431_ heichips25_sap3/_1036_ heichips25_sap3/_1018_ heichips25_sap3/_1037_
+ VPWR VGND sg13g2_xor2_1
Xheichips25_sap3__3362_ heichips25_sap3/_0971_ heichips25_sap3/_0967_ heichips25_sap3/_0970_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__2313_ heichips25_sap3/_1713_ heichips25_sap3/_1732_ heichips25_sap3/_1695_
+ heichips25_sap3/_1734_ VPWR VGND sg13g2_nand3_1
XFILLER_44_742 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3293_ VGND VPWR heichips25_sap3/net127 heichips25_sap3/_0901_ heichips25_sap3/_0905_
+ heichips25_sap3/_0904_ sg13g2_a21oi_1
Xheichips25_sap3__2244_ heichips25_sap3/_1665_ heichips25_sap3/_1559_ heichips25_sap3/_1664_
+ VPWR VGND sg13g2_nand2_1
XFILLER_44_786 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2175_ VPWR heichips25_sap3/_1596_ heichips25_sap3/_1595_ VGND sg13g2_inv_1
XFILLER_31_403 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__1959_ VPWR heichips25_sap3/_1385_ heichips25_sap3__3932_/Q VGND
+ sg13g2_inv_1
Xheichips25_can_lehmann_fsm__2855__786 VPWR VGND net785 sg13g2_tiehi
XFILLER_3_392 VPWR VGND sg13g2_fill_1
XFILLER_26_1021 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3629_ heichips25_sap3/_0127_ heichips25_sap3/_1130_ heichips25_sap3/_1186_
+ heichips25_sap3/net103 heichips25_sap3/_1423_ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2850_ net795 VGND VPWR heichips25_can_lehmann_fsm/_0075_
+ heichips25_can_lehmann_fsm__2850_/Q clknet_leaf_8_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2781_ net644 VGND VPWR heichips25_can_lehmann_fsm/net1261
+ heichips25_can_lehmann_fsm__2781_/Q clknet_leaf_4_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1801_ heichips25_can_lehmann_fsm/net338 heichips25_can_lehmann_fsm/_0989_
+ heichips25_can_lehmann_fsm__2900_/Q heichips25_can_lehmann_fsm/_1117_ VPWR VGND
+ sg13g2_nand3_1
Xheichips25_can_lehmann_fsm__1732_ heichips25_can_lehmann_fsm__2833_/Q heichips25_can_lehmann_fsm__2832_/Q
+ heichips25_can_lehmann_fsm__2831_/Q heichips25_can_lehmann_fsm__2830_/Q heichips25_can_lehmann_fsm/_1053_
+ VPWR VGND sg13g2_nor4_1
XFILLER_34_241 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1663_ VPWR heichips25_can_lehmann_fsm/_0987_ net5 VGND
+ sg13g2_inv_1
Xheichips25_can_lehmann_fsm__1594_ VPWR heichips25_can_lehmann_fsm/_0918_ heichips25_can_lehmann_fsm/net863
+ VGND sg13g2_inv_1
XFILLER_23_959 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2215_ heichips25_can_lehmann_fsm/net329 VPWR heichips25_can_lehmann_fsm/_0543_
+ VGND heichips25_can_lehmann_fsm/net1186 heichips25_can_lehmann_fsm/net162 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2146_ heichips25_can_lehmann_fsm/_0485_ heichips25_can_lehmann_fsm/net337
+ heichips25_can_lehmann_fsm/_0483_ heichips25_can_lehmann_fsm/net316 heichips25_can_lehmann_fsm__2926_/Q
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2077_ heichips25_can_lehmann_fsm/net322 VPWR heichips25_can_lehmann_fsm/_0422_
+ VGND heichips25_can_lehmann_fsm/net346 heichips25_can_lehmann_fsm/net179 sg13g2_o21ai_1
XFILLER_45_517 VPWR VGND sg13g2_fill_2
XFILLER_45_506 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2979_ net708 VGND VPWR heichips25_can_lehmann_fsm/_0204_
+ heichips25_can_lehmann_fsm__2979_/Q clknet_leaf_12_clk sg13g2_dfrbpq_1
Xheichips25_sap3_fanout141 heichips25_sap3/net143 heichips25_sap3/net141 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout130 heichips25_sap3/_0719_ heichips25_sap3/net130 VPWR VGND
+ sg13g2_buf_1
XFILLER_43_11 VPWR VGND sg13g2_decap_8
Xheichips25_sap3_fanout152 heichips25_sap3/_0718_ heichips25_sap3/net152 VPWR VGND
+ sg13g2_buf_1
XFILLER_25_274 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm_hold1220 heichips25_can_lehmann_fsm__2796_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1219 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1231 heichips25_can_lehmann_fsm/_0269_ VPWR VGND heichips25_can_lehmann_fsm/net1230
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1242 heichips25_can_lehmann_fsm/_0012_ VPWR VGND heichips25_can_lehmann_fsm/net1241
+ sg13g2_dlygate4sd3_1
XFILLER_43_99 VPWR VGND sg13g2_fill_2
XFILLER_41_778 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_hold1275 heichips25_can_lehmann_fsm__2794_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1274 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1264 heichips25_can_lehmann_fsm/_0003_ VPWR VGND heichips25_can_lehmann_fsm/net1263
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1253 heichips25_can_lehmann_fsm/_0010_ VPWR VGND heichips25_can_lehmann_fsm/net1252
+ sg13g2_dlygate4sd3_1
XFILLER_9_429 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3980_ heichips25_sap3/net434 VGND VPWR heichips25_sap3/_0121_ heichips25_sap3__3980_/Q
+ heichips25_sap3__4012_/CLK sg13g2_dfrbpq_1
Xheichips25_sap3__2931_ heichips25_sap3/_0567_ heichips25_sap3/_0568_ heichips25_sap3/_0566_
+ heichips25_sap3/_0570_ VPWR VGND heichips25_sap3/_0569_ sg13g2_nand4_1
Xheichips25_sap3__2862_ heichips25_sap3/_1367_ VPWR heichips25_sap3/_0504_ VGND heichips25_sap3/_1619_
+ heichips25_sap3/_1714_ sg13g2_o21ai_1
XFILLER_4_123 VPWR VGND sg13g2_decap_8
XFILLER_49_1010 VPWR VGND sg13g2_decap_8
XFILLER_4_167 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2793_ heichips25_sap3/_1721_ heichips25_sap3/_1886_ heichips25_sap3/_0438_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__3414_ heichips25_sap3/_1021_ heichips25_sap3/_1020_ heichips25_sap3/_0873_
+ VPWR VGND sg13g2_nand2b_1
XFILLER_36_517 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3345_ uio_oe_sap3\[3\] heichips25_sap3/_0884_ heichips25_sap3/_0955_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__3276_ heichips25_sap3/_0889_ heichips25_sap3/_0732_ heichips25_sap3/net166
+ VPWR VGND sg13g2_nand2_1
XFILLER_44_583 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2227_ heichips25_sap3/_1639_ heichips25_sap3/net220 heichips25_sap3/_1647_
+ heichips25_sap3/_1648_ VPWR VGND sg13g2_nor3_1
XFILLER_17_786 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2158_ heichips25_sap3/_1577_ heichips25_sap3/_1578_ heichips25_sap3/_1579_
+ VPWR VGND sg13g2_nor2_1
XFILLER_31_255 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2089_ heichips25_sap3/_1505_ heichips25_sap3/_1507_ heichips25_sap3/_1445_
+ heichips25_sap3/_1510_ VPWR VGND sg13g2_nand3_1
XFILLER_31_288 VPWR VGND sg13g2_decap_8
XFILLER_8_451 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2000_ heichips25_can_lehmann_fsm/net326 VPWR heichips25_can_lehmann_fsm/_0356_
+ VGND heichips25_can_lehmann_fsm/net1251 heichips25_can_lehmann_fsm/net180 sg13g2_o21ai_1
XFILLER_4_690 VPWR VGND sg13g2_fill_1
XFILLER_39_344 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2902_ net691 VGND VPWR heichips25_can_lehmann_fsm/_0127_
+ heichips25_can_lehmann_fsm__2902_/Q clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_39_366 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2833_ net540 VGND VPWR heichips25_can_lehmann_fsm/_0058_
+ heichips25_can_lehmann_fsm__2833_/Q clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_27_539 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2764_ heichips25_can_lehmann_fsm/net487 VPWR heichips25_can_lehmann_fsm/_0848_
+ VGND heichips25_can_lehmann_fsm/net1116 heichips25_can_lehmann_fsm/net378 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__1715_ heichips25_can_lehmann_fsm/_1038_ VPWR uo_out_fsm\[0\]
+ VGND heichips25_can_lehmann_fsm/_0977_ heichips25_can_lehmann_fsm/_1033_ sg13g2_o21ai_1
XFILLER_23_701 VPWR VGND sg13g2_fill_2
XFILLER_23_712 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2695_ VGND VPWR heichips25_can_lehmann_fsm/_0872_ heichips25_can_lehmann_fsm/net404
+ heichips25_can_lehmann_fsm/_0247_ heichips25_can_lehmann_fsm/_0813_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__1646_ VPWR heichips25_can_lehmann_fsm/_0970_ heichips25_can_lehmann_fsm/net895
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__1577_ VPWR heichips25_can_lehmann_fsm/_0901_ heichips25_can_lehmann_fsm/net885
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__2129_ heichips25_can_lehmann_fsm/_1090_ VPWR heichips25_can_lehmann_fsm/_0468_
+ VGND heichips25_can_lehmann_fsm/net219 heichips25_can_lehmann_fsm/_0467_ sg13g2_o21ai_1
XFILLER_45_347 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3130_ heichips25_sap3/_0643_ heichips25_sap3/_0742_ heichips25_sap3/_0743_
+ VPWR VGND sg13g2_and2_1
Xheichips25_sap3__3061_ heichips25_sap3/_0674_ heichips25_sap3/_1605_ heichips25_sap3/_1664_
+ heichips25_sap3/_1517_ heichips25_sap3/_1496_ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2984__689 VPWR VGND net688 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__3045__679 VPWR VGND net678 sg13g2_tiehi
XFILLER_41_520 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2012_ heichips25_sap3/net1019 heichips25_sap3/net342 heichips25_sap3__4058_/Q
+ heichips25_sap3/_0017_ VPWR VGND heichips25_sap3__4047_/Q sg13g2_nand4_1
XFILLER_13_222 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm_hold1050 heichips25_can_lehmann_fsm__2913_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1049 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1083 heichips25_can_lehmann_fsm__2952_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1082 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1061 heichips25_can_lehmann_fsm__2949_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1060 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1094 heichips25_can_lehmann_fsm__2835_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1093 sg13g2_dlygate4sd3_1
XFILLER_10_940 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3963_ heichips25_sap3/net443 VGND VPWR heichips25_sap3/_0104_ heichips25_sap3__3963_/Q
+ clkload19/A sg13g2_dfrbpq_1
Xclkload29 VPWR clkload29/Y clkload29/A VGND sg13g2_inv_1
XFILLER_5_421 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2914_ heichips25_sap3/_0554_ heichips25_sap3/_1382_ heichips25_sap3/net211
+ VPWR VGND sg13g2_xnor2_1
Xclkload18 VPWR clkload18/Y clkload18/A VGND sg13g2_inv_1
Xheichips25_sap3__3894_ heichips25_sap3/net448 VGND VPWR heichips25_sap3/_0035_ heichips25_sap3__3894_/Q
+ net818 sg13g2_dfrbpq_1
Xheichips25_sap3__2845_ VGND VPWR heichips25_sap3/net154 heichips25_sap3/_0403_ heichips25_sap3/_0488_
+ heichips25_sap3/_0487_ sg13g2_a21oi_1
Xheichips25_sap3__2776_ heichips25_sap3/_0418_ heichips25_sap3/_0419_ heichips25_sap3/_0384_
+ heichips25_sap3/_0422_ VPWR VGND heichips25_sap3/_0421_ sg13g2_nand4_1
XFILLER_1_671 VPWR VGND sg13g2_fill_1
XFILLER_0_192 VPWR VGND sg13g2_decap_8
XFILLER_48_163 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3328_ heichips25_sap3/_0938_ heichips25_sap3__3942_/Q heichips25_sap3/net105
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__3259_ heichips25_sap3/net61 heichips25_sap3/_0867_ heichips25_sap3/_0872_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_can_lehmann_fsm__2480_ heichips25_can_lehmann_fsm/net482 VPWR heichips25_can_lehmann_fsm/_0706_
+ VGND heichips25_can_lehmann_fsm/net869 heichips25_can_lehmann_fsm/net370 sg13g2_o21ai_1
XFILLER_9_760 VPWR VGND sg13g2_fill_1
XFILLER_8_292 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__3032_ net597 VGND VPWR heichips25_can_lehmann_fsm/_0257_
+ heichips25_can_lehmann_fsm__3032_/Q clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_27_325 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2816_ net574 VGND VPWR heichips25_can_lehmann_fsm/net1222
+ heichips25_can_lehmann_fsm__2816_/Q clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_27_347 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2747_ VGND VPWR heichips25_can_lehmann_fsm/_0858_ heichips25_can_lehmann_fsm/net421
+ heichips25_can_lehmann_fsm/_0273_ heichips25_can_lehmann_fsm/_0839_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm_hold925 heichips25_can_lehmann_fsm__3014_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net924 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__2678_ heichips25_can_lehmann_fsm/net464 VPWR heichips25_can_lehmann_fsm/_0805_
+ VGND heichips25_can_lehmann_fsm/net924 heichips25_can_lehmann_fsm/net394 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm_hold903 heichips25_can_lehmann_fsm__2966_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net902 sg13g2_dlygate4sd3_1
XFILLER_11_715 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm_hold914 heichips25_can_lehmann_fsm__2897_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net913 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__1629_ VPWR heichips25_can_lehmann_fsm/_0953_ heichips25_can_lehmann_fsm/net1167
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm_hold936 heichips25_can_lehmann_fsm/_0172_ VPWR VGND heichips25_can_lehmann_fsm/net935
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold947 heichips25_can_lehmann_fsm__2971_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net946 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold958 heichips25_can_lehmann_fsm__2973_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net957 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold969 heichips25_can_lehmann_fsm__2858_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net968 sg13g2_dlygate4sd3_1
XFILLER_6_207 VPWR VGND sg13g2_decap_8
XFILLER_10_269 VPWR VGND sg13g2_decap_8
XFILLER_6_4 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2630_ heichips25_sap3/_1487_ heichips25_sap3/_1502_ heichips25_sap3/net237
+ heichips25_sap3/_0297_ VPWR VGND heichips25_sap3/_1541_ sg13g2_nand4_1
XFILLER_2_457 VPWR VGND sg13g2_decap_4
XFILLER_49_32 VPWR VGND sg13g2_decap_8
XFILLER_2_479 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2561_ heichips25_sap3/_0236_ heichips25_sap3/net75 heichips25_sap3__3990_/Q
+ heichips25_sap3/net216 heichips25_sap3__4014_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2492_ VGND VPWR heichips25_sap3__3940_/Q heichips25_sap3/net88 heichips25_sap3/_1905_
+ heichips25_sap3/net89 sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2949__540 VPWR VGND net539 sg13g2_tiehi
XFILLER_45_144 VPWR VGND sg13g2_fill_1
XFILLER_18_358 VPWR VGND sg13g2_fill_1
XFILLER_46_678 VPWR VGND sg13g2_decap_4
XFILLER_45_177 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3113_ heichips25_sap3/_1509_ VPWR heichips25_sap3/_0726_ VGND heichips25_sap3/net230
+ heichips25_sap3/_1607_ sg13g2_o21ai_1
XFILLER_33_306 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3044_ heichips25_sap3/net263 VPWR heichips25_sap3/_0657_ VGND heichips25_sap3/_0654_
+ heichips25_sap3/_0655_ sg13g2_o21ai_1
XFILLER_14_542 VPWR VGND sg13g2_decap_8
XFILLER_10_781 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3946_ heichips25_sap3/net444 VGND VPWR heichips25_sap3/_0087_ heichips25_sap3__3946_/Q
+ heichips25_sap3__4024_/CLK sg13g2_dfrbpq_1
XFILLER_5_240 VPWR VGND sg13g2_decap_8
XFILLER_6_785 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2828_ VGND VPWR heichips25_sap3/net64 heichips25_sap3/_0468_ heichips25_sap3/_0472_
+ heichips25_sap3/net204 sg13g2_a21oi_1
Xheichips25_sap3__2759_ heichips25_sap3/_0361_ heichips25_sap3/_0377_ heichips25_sap3/_0402_
+ heichips25_sap3/_0405_ VPWR VGND sg13g2_nor3_1
Xheichips25_can_lehmann_fsm__1980_ VPWR VGND heichips25_can_lehmann_fsm/net196 heichips25_can_lehmann_fsm/_0338_
+ heichips25_can_lehmann_fsm/_0337_ heichips25_can_lehmann_fsm/_0333_ heichips25_can_lehmann_fsm/_0007_
+ heichips25_can_lehmann_fsm/_0336_ sg13g2_a221oi_1
XFILLER_49_483 VPWR VGND sg13g2_decap_4
Xinput5 ui_in[2] net5 VPWR VGND sg13g2_buf_1
XFILLER_25_807 VPWR VGND sg13g2_fill_1
XFILLER_36_155 VPWR VGND sg13g2_decap_4
XFILLER_24_306 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2928__624 VPWR VGND net623 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2601_ VGND VPWR heichips25_can_lehmann_fsm/_0897_ heichips25_can_lehmann_fsm/net366
+ heichips25_can_lehmann_fsm/_0200_ heichips25_can_lehmann_fsm/_0766_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2532_ heichips25_can_lehmann_fsm/net477 VPWR heichips25_can_lehmann_fsm/_0732_
+ VGND heichips25_can_lehmann_fsm/net1005 heichips25_can_lehmann_fsm/net368 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2463_ VGND VPWR heichips25_can_lehmann_fsm/_0932_ heichips25_can_lehmann_fsm/net422
+ heichips25_can_lehmann_fsm/_0131_ heichips25_can_lehmann_fsm/_0697_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2394_ heichips25_can_lehmann_fsm/net470 VPWR heichips25_can_lehmann_fsm/_0663_
+ VGND heichips25_can_lehmann_fsm/net1066 heichips25_can_lehmann_fsm/net390 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__3015_ net762 VGND VPWR heichips25_can_lehmann_fsm/_0240_
+ heichips25_can_lehmann_fsm__3015_/Q clknet_leaf_19_clk sg13g2_dfrbpq_1
XFILLER_47_409 VPWR VGND sg13g2_fill_2
XFILLER_19_46 VPWR VGND sg13g2_fill_2
XFILLER_28_601 VPWR VGND sg13g2_fill_2
XFILLER_28_612 VPWR VGND sg13g2_decap_8
XFILLER_28_634 VPWR VGND sg13g2_decap_8
XFILLER_43_626 VPWR VGND sg13g2_fill_1
XFILLER_16_829 VPWR VGND sg13g2_fill_1
XFILLER_15_328 VPWR VGND sg13g2_fill_2
XFILLER_27_199 VPWR VGND sg13g2_fill_1
XFILLER_30_309 VPWR VGND sg13g2_fill_2
XFILLER_11_545 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__1992_ VPWR heichips25_sap3/_1418_ heichips25_sap3__3953_/Q VGND
+ sg13g2_inv_1
Xheichips25_sap3__3800_ VPWR VGND heichips25_sap3__3942_/Q heichips25_sap3/_1308_
+ heichips25_sap3/_1274_ heichips25_sap3__3982_/Q heichips25_sap3/_1309_ heichips25_sap3/_1259_
+ sg13g2_a221oi_1
Xheichips25_sap3__3731_ heichips25_sap3__4030_/Q heichips25_sap3/net1031 heichips25_sap3/_1248_
+ VPWR VGND heichips25_sap3__4029_/Q sg13g2_nand3b_1
Xclkbuf_4_14_0_heichips25_sap3\_sap_3_inst.alu_inst.clk clknet_0_heichips25_sap3\/sap_3_inst.alu_inst.clk
+ clknet_4_14_0_heichips25_sap3\/sap_3_inst.alu_inst.clk VPWR VGND sg13g2_buf_8
XFILLER_3_722 VPWR VGND sg13g2_decap_8
XFILLER_2_221 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3662_ uio_oe_sap3\[3\] heichips25_sap3/net112 heichips25_sap3/_1207_
+ heichips25_sap3/_1208_ VPWR VGND sg13g2_nor3_1
Xheichips25_sap3__3593_ heichips25_sap3/net101 heichips25_sap3/_1167_ heichips25_sap3/_1168_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__2613_ heichips25_sap3/_1484_ heichips25_sap3/_1579_ heichips25_sap3/net241
+ heichips25_sap3/_0284_ VPWR VGND heichips25_sap3/_1612_ sg13g2_nand4_1
Xheichips25_sap3__2544_ heichips25_sap3/_0218_ heichips25_sap3/_0219_ heichips25_sap3/_0214_
+ heichips25_sap3/_0220_ VPWR VGND sg13g2_nand3_1
XFILLER_47_932 VPWR VGND sg13g2_fill_2
XFILLER_47_976 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2475_ heichips25_sap3/_1888_ heichips25_sap3__3927_/Q heichips25_sap3/_1881_
+ VPWR VGND sg13g2_nand2_1
XFILLER_18_111 VPWR VGND sg13g2_fill_1
XFILLER_47_987 VPWR VGND sg13g2_fill_2
XFILLER_47_998 VPWR VGND sg13g2_fill_1
XFILLER_19_689 VPWR VGND sg13g2_fill_1
XFILLER_33_114 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3027_ heichips25_sap3/_1525_ heichips25_sap3/_1535_ heichips25_sap3/_0639_
+ heichips25_sap3/_0640_ VPWR VGND sg13g2_nor3_1
XFILLER_30_876 VPWR VGND sg13g2_decap_4
XFILLER_6_560 VPWR VGND sg13g2_decap_4
XFILLER_6_593 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3929_ heichips25_sap3/net435 VGND VPWR heichips25_sap3/_0070_ heichips25_sap3__3929_/Q
+ clkload23/A sg13g2_dfrbpq_1
Xheichips25_sap3_clk_div_param_inst__1_ VPWR heichips25_sap3_clk_div_param_inst__2_/D
+ heichips25_sap3_clk_div_param_inst__1_/A VGND sg13g2_inv_1
XFILLER_2_60 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1963_ heichips25_can_lehmann_fsm__2797_/Q heichips25_can_lehmann_fsm/net181
+ heichips25_can_lehmann_fsm/_0324_ VPWR VGND sg13g2_nor2_1
Xheichips25_can_lehmann_fsm__1894_ heichips25_can_lehmann_fsm/_1207_ heichips25_can_lehmann_fsm/_0896_
+ heichips25_can_lehmann_fsm/net349 VPWR VGND sg13g2_nand2_1
Xheichips25_can_lehmann_fsm__2865__766 VPWR VGND net765 sg13g2_tiehi
Xheichips25_sap3_hold1126 heichips25_sap3/_0195_ VPWR VGND heichips25_sap3/net1125
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__2515_ VGND VPWR heichips25_can_lehmann_fsm/_0919_ heichips25_can_lehmann_fsm/net426
+ heichips25_can_lehmann_fsm/_0157_ heichips25_can_lehmann_fsm/_0723_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2446_ heichips25_can_lehmann_fsm/net468 VPWR heichips25_can_lehmann_fsm/_0689_
+ VGND heichips25_can_lehmann_fsm__2898_/Q heichips25_can_lehmann_fsm/net398 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2377_ VGND VPWR heichips25_can_lehmann_fsm/_0957_ heichips25_can_lehmann_fsm/net383
+ heichips25_can_lehmann_fsm/_0088_ heichips25_can_lehmann_fsm/_0654_ sg13g2_a21oi_1
XFILLER_20_397 VPWR VGND sg13g2_fill_1
XFILLER_21_25 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm_fanout430 heichips25_can_lehmann_fsm/net431 heichips25_can_lehmann_fsm/net430
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout474 heichips25_can_lehmann_fsm/net475 heichips25_can_lehmann_fsm/net474
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout496 heichips25_can_lehmann_fsm/net503 heichips25_can_lehmann_fsm/net496
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout485 heichips25_can_lehmann_fsm/net489 heichips25_can_lehmann_fsm/net485
+ VPWR VGND sg13g2_buf_1
XFILLER_47_217 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2260_ heichips25_sap3/_1681_ heichips25_sap3/_1551_ heichips25_sap3/net246
+ heichips25_sap3/_1546_ heichips25_sap3/_1459_ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2191_ heichips25_sap3/_1612_ heichips25_sap3/_1500_ heichips25_sap3/_1513_
+ VPWR VGND sg13g2_nand2_1
XFILLER_28_497 VPWR VGND sg13g2_fill_2
XFILLER_24_670 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__1975_ VPWR heichips25_sap3/_1401_ heichips25_sap3__4015_/Q VGND
+ sg13g2_inv_1
Xheichips25_sap3__3714_ heichips25_sap3/_0158_ heichips25_sap3/_1124_ heichips25_sap3/_1240_
+ heichips25_sap3/net114 heichips25_sap3/_1413_ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3645_ heichips25_sap3/_1083_ heichips25_sap3__3994_/Q heichips25_sap3/_1187_
+ heichips25_sap3/_0135_ VPWR VGND sg13g2_mux2_1
XFILLER_3_585 VPWR VGND sg13g2_decap_4
XFILLER_3_574 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3576_ heichips25_sap3/net100 heichips25_sap3/_0924_ heichips25_sap3/_1154_
+ heichips25_sap3/_1155_ VPWR VGND sg13g2_nor3_1
XFILLER_47_751 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2527_ heichips25_sap3/_0204_ heichips25_sap3/net78 heichips25_sap3__4019_/Q
+ heichips25_sap3/net89 heichips25_sap3__3939_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2458_ heichips25_sap3/net230 heichips25_sap3/_1559_ heichips25_sap3/_1871_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__2389_ heichips25_sap3/_1808_ heichips25_sap3/_1806_ heichips25_sap3/_1807_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__4059_ heichips25_sap3/net453 VGND VPWR heichips25_sap3__4059_/D
+ heichips25_sap3__4059_/Q clknet_leaf_22_clk sg13g2_dfrbpq_1
XFILLER_15_692 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2300_ VGND VPWR heichips25_can_lehmann_fsm/_0607_ heichips25_can_lehmann_fsm/net1201
+ heichips25_can_lehmann_fsm/_0055_ heichips25_can_lehmann_fsm/_0610_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2231_ heichips25_can_lehmann_fsm/_0555_ heichips25_can_lehmann_fsm/_0496_
+ heichips25_can_lehmann_fsm/_0554_ heichips25_can_lehmann_fsm/net176 heichips25_can_lehmann_fsm/net1002
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2162_ heichips25_can_lehmann_fsm/_0501_ heichips25_can_lehmann_fsm/net164
+ heichips25_can_lehmann_fsm/_0975_ heichips25_can_lehmann_fsm/net175 heichips25_can_lehmann_fsm/net1204
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2093_ VGND VPWR net16 heichips25_can_lehmann_fsm/net195
+ heichips25_can_lehmann_fsm/_0435_ heichips25_can_lehmann_fsm/net182 sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2995_ net633 VGND VPWR heichips25_can_lehmann_fsm/net929
+ heichips25_can_lehmann_fsm__2995_/Q clknet_leaf_21_clk sg13g2_dfrbpq_1
XFILLER_38_751 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1946_ heichips25_can_lehmann_fsm/_0309_ heichips25_can_lehmann_fsm/_1215_
+ heichips25_can_lehmann_fsm/_1234_ heichips25_can_lehmann_fsm/_0303_ VPWR VGND sg13g2_and3_1
Xheichips25_can_lehmann_fsm__3043__711 VPWR VGND net710 sg13g2_tiehi
XFILLER_26_946 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1877_ heichips25_can_lehmann_fsm/_1191_ heichips25_can_lehmann_fsm/net295
+ heichips25_can_lehmann_fsm__2964_/Q heichips25_can_lehmann_fsm/net332 heichips25_can_lehmann_fsm__3036_/Q
+ VPWR VGND sg13g2_a22oi_1
XFILLER_16_69 VPWR VGND sg13g2_fill_2
XFILLER_5_806 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2429_ VGND VPWR heichips25_can_lehmann_fsm/_0940_ heichips25_can_lehmann_fsm/net372
+ heichips25_can_lehmann_fsm/_0114_ heichips25_can_lehmann_fsm/_0680_ sg13g2_a21oi_1
XFILLER_4_338 VPWR VGND sg13g2_fill_2
XFILLER_0_522 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3430_ heichips25_sap3/_1036_ heichips25_sap3/_1030_ heichips25_sap3/_1035_
+ heichips25_sap3/net125 heichips25_sap3/_1420_ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3361_ heichips25_sap3/_0970_ heichips25_sap3/net59 heichips25_sap3/_0969_
+ VPWR VGND sg13g2_nand2b_1
Xheichips25_sap3__2312_ heichips25_sap3/_1680_ heichips25_sap3/_1693_ heichips25_sap3/_1712_
+ heichips25_sap3/_1731_ heichips25_sap3/_1733_ VPWR VGND sg13g2_nor4_1
Xheichips25_sap3__3292_ heichips25_sap3/net127 heichips25_sap3/_0903_ heichips25_sap3/_0904_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__2243_ VGND VPWR heichips25_sap3/_1664_ heichips25_sap3/_1557_ heichips25_sap3/_1522_
+ sg13g2_or2_1
XFILLER_28_261 VPWR VGND sg13g2_fill_2
XFILLER_43_286 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2174_ VGND VPWR heichips25_sap3/_1504_ heichips25_sap3/_1525_ heichips25_sap3/_1595_
+ heichips25_sap3/_1570_ sg13g2_a21oi_1
XFILLER_8_600 VPWR VGND sg13g2_decap_4
XFILLER_11_161 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2959__789 VPWR VGND net788 sg13g2_tiehi
Xheichips25_sap3__1958_ VPWR heichips25_sap3/_1384_ heichips25_sap3/net276 VGND sg13g2_inv_1
Xheichips25_sap3__3628_ heichips25_sap3/net142 heichips25_sap3/_1082_ heichips25_sap3/_1186_
+ VPWR VGND sg13g2_and2_1
XFILLER_21_4 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3559_ heichips25_sap3__3961_/Q heichips25_sap3/_1141_ heichips25_sap3/_1134_
+ heichips25_sap3/_0102_ VPWR VGND sg13g2_mux2_1
Xheichips25_can_lehmann_fsm__2780_ net646 VGND VPWR heichips25_can_lehmann_fsm/net1250
+ heichips25_can_lehmann_fsm__2780_/Q clknet_leaf_2_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1800_ VPWR VGND heichips25_can_lehmann_fsm__2948_/Q heichips25_can_lehmann_fsm/_1115_
+ heichips25_can_lehmann_fsm/net306 heichips25_can_lehmann_fsm__3020_/Q heichips25_can_lehmann_fsm/_1116_
+ heichips25_can_lehmann_fsm/net310 sg13g2_a221oi_1
XFILLER_47_581 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1731_ heichips25_can_lehmann_fsm/net1158 heichips25_can_lehmann_fsm__2830_/Q
+ heichips25_can_lehmann_fsm/_1051_ heichips25_can_lehmann_fsm/_1052_ VPWR VGND sg13g2_nor3_1
XFILLER_23_949 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1662_ VPWR heichips25_can_lehmann_fsm/_0986_ net4 VGND
+ sg13g2_inv_1
XFILLER_34_264 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1593_ VPWR heichips25_can_lehmann_fsm/_0917_ heichips25_can_lehmann_fsm/net1106
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__2214_ heichips25_can_lehmann_fsm/_0542_ heichips25_can_lehmann_fsm/net165
+ heichips25_can_lehmann_fsm/_0541_ heichips25_can_lehmann_fsm/net176 heichips25_can_lehmann_fsm/net1006
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2145_ heichips25_can_lehmann_fsm/_0484_ heichips25_can_lehmann_fsm/net334
+ heichips25_can_lehmann_fsm__3046_/Q heichips25_can_lehmann_fsm/net299 heichips25_can_lehmann_fsm__2902_/Q
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2076_ heichips25_can_lehmann_fsm/_0421_ heichips25_can_lehmann_fsm/net186
+ heichips25_can_lehmann_fsm/_0420_ heichips25_can_lehmann_fsm/net195 net13 VPWR VGND
+ sg13g2_a22oi_1
XFILLER_38_570 VPWR VGND sg13g2_decap_8
XFILLER_26_721 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2978_ net712 VGND VPWR heichips25_can_lehmann_fsm/_0203_
+ heichips25_can_lehmann_fsm__2978_/Q clknet_leaf_13_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1929_ heichips25_can_lehmann_fsm/_0291_ VPWR heichips25_can_lehmann_fsm/_0292_
+ VGND heichips25_can_lehmann_fsm__2888_/Q heichips25_can_lehmann_fsm/net336 sg13g2_o21ai_1
Xheichips25_sap3_fanout131 heichips25_sap3/_0881_ heichips25_sap3/net131 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout120 heichips25_sap3/_0750_ heichips25_sap3/net120 VPWR VGND
+ sg13g2_buf_1
XFILLER_41_724 VPWR VGND sg13g2_fill_2
Xheichips25_sap3_fanout142 heichips25_sap3/net143 heichips25_sap3/net142 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout153 heichips25_sap3/_0606_ heichips25_sap3/net153 VPWR VGND
+ sg13g2_buf_1
XFILLER_14_949 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_hold1232 heichips25_can_lehmann_fsm__2814_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1231 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1221 heichips25_can_lehmann_fsm/_0022_ VPWR VGND heichips25_can_lehmann_fsm/net1220
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1210 heichips25_can_lehmann_fsm__2828_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1209 sg13g2_dlygate4sd3_1
XFILLER_13_437 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm_hold1265 heichips25_can_lehmann_fsm__2798_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1264 sg13g2_dlygate4sd3_1
XFILLER_43_78 VPWR VGND sg13g2_fill_1
XFILLER_40_245 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_hold1243 heichips25_can_lehmann_fsm__2778_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1242 sg13g2_dlygate4sd3_1
XFILLER_22_960 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm_hold1254 heichips25_can_lehmann_fsm__2779_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1253 sg13g2_dlygate4sd3_1
XFILLER_22_993 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2930_ heichips25_sap3/net159 VPWR heichips25_sap3/_0569_ VGND heichips25_sap3/net276
+ heichips25_sap3__3921_/Q sg13g2_o21ai_1
Xheichips25_sap3__2861_ heichips25_sap3/_0482_ VPWR heichips25_sap3/_0503_ VGND heichips25_sap3/_0483_
+ heichips25_sap3/_0484_ sg13g2_o21ai_1
Xheichips25_sap3__2792_ heichips25_sap3/_1877_ heichips25_sap3/net158 heichips25_sap3/net204
+ heichips25_sap3/_0437_ VPWR VGND sg13g2_nor3_1
XFILLER_49_802 VPWR VGND sg13g2_fill_2
XFILLER_48_301 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3413_ heichips25_sap3/_0794_ VPWR heichips25_sap3/_1020_ VGND heichips25_sap3/net62
+ heichips25_sap3/_0868_ sg13g2_o21ai_1
XFILLER_1_1024 VPWR VGND sg13g2_decap_4
XFILLER_29_570 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3344_ VGND VPWR heichips25_sap3/_0952_ heichips25_sap3/_0953_ heichips25_sap3/_0954_
+ heichips25_sap3/net120 sg13g2_a21oi_1
Xheichips25_sap3__3275_ heichips25_sap3/_0731_ heichips25_sap3/net166 heichips25_sap3/_0888_
+ VPWR VGND sg13g2_nor2b_1
XFILLER_44_562 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2226_ VGND VPWR heichips25_sap3/net237 heichips25_sap3/_1620_ heichips25_sap3/_1647_
+ heichips25_sap3/_1646_ sg13g2_a21oi_1
XFILLER_16_275 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2157_ heichips25_sap3/net234 heichips25_sap3/_1475_ heichips25_sap3/_1578_
+ VPWR VGND sg13g2_nor2_1
XFILLER_16_297 VPWR VGND sg13g2_fill_2
XFILLER_31_234 VPWR VGND sg13g2_decap_8
XFILLER_8_430 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2088_ heichips25_sap3/_1446_ heichips25_sap3/_1506_ heichips25_sap3/_1508_
+ heichips25_sap3/_1509_ VPWR VGND sg13g2_nor3_1
XFILLER_31_278 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2901_ net693 VGND VPWR heichips25_can_lehmann_fsm/net1009
+ heichips25_can_lehmann_fsm__2901_/Q clknet_leaf_6_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2832_ net542 VGND VPWR heichips25_can_lehmann_fsm/net1190
+ heichips25_can_lehmann_fsm__2832_/Q clknet_leaf_9_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2763_ VGND VPWR heichips25_can_lehmann_fsm/_0854_ heichips25_can_lehmann_fsm/net417
+ heichips25_can_lehmann_fsm/_0281_ heichips25_can_lehmann_fsm/_0847_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2694_ heichips25_can_lehmann_fsm/net472 VPWR heichips25_can_lehmann_fsm/_0813_
+ VGND heichips25_can_lehmann_fsm/net849 heichips25_can_lehmann_fsm/net404 sg13g2_o21ai_1
XFILLER_35_573 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__1714_ VGND VPWR heichips25_can_lehmann_fsm__2785_/Q heichips25_can_lehmann_fsm/_1037_
+ heichips25_can_lehmann_fsm/_1038_ heichips25_can_lehmann_fsm/_1036_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__1645_ VPWR heichips25_can_lehmann_fsm/_0969_ heichips25_can_lehmann_fsm/net1099
+ VGND sg13g2_inv_1
XFILLER_22_223 VPWR VGND sg13g2_fill_2
XFILLER_22_256 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1576_ VPWR heichips25_can_lehmann_fsm/_0900_ heichips25_can_lehmann_fsm/net887
+ VGND sg13g2_inv_1
XFILLER_13_59 VPWR VGND sg13g2_decap_4
XFILLER_2_606 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2128_ heichips25_can_lehmann_fsm/_0466_ VPWR heichips25_can_lehmann_fsm/_0467_
+ VGND heichips25_can_lehmann_fsm__2880_/Q heichips25_can_lehmann_fsm/net335 sg13g2_o21ai_1
XFILLER_49_109 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2059_ heichips25_can_lehmann_fsm/_0407_ heichips25_can_lehmann_fsm/net196
+ heichips25_can_lehmann_fsm/_0406_ heichips25_can_lehmann_fsm/net200 heichips25_can_lehmann_fsm__2801_/Q
+ VPWR VGND sg13g2_a22oi_1
XFILLER_38_56 VPWR VGND sg13g2_decap_8
XFILLER_46_838 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3060_ heichips25_sap3/_0673_ heichips25_sap3/net266 heichips25_sap3/_1773_
+ VPWR VGND sg13g2_nand2_1
XFILLER_26_562 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2011_ heichips25_sap3/_1433_ heichips25_sap3/net342 heichips25_sap3/net1138
+ VPWR VGND sg13g2_nand2_1
XFILLER_13_201 VPWR VGND sg13g2_decap_8
XFILLER_26_595 VPWR VGND sg13g2_decap_4
XFILLER_13_245 VPWR VGND sg13g2_decap_4
XFILLER_13_256 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm_hold1040 heichips25_can_lehmann_fsm__3031_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1039 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1051 heichips25_can_lehmann_fsm__2847_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1050 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1062 heichips25_can_lehmann_fsm/_0175_ VPWR VGND heichips25_can_lehmann_fsm/net1061
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1084 heichips25_can_lehmann_fsm__2963_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1083 sg13g2_dlygate4sd3_1
XFILLER_9_227 VPWR VGND sg13g2_decap_4
XFILLER_16_1021 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3962_ heichips25_sap3/net444 VGND VPWR heichips25_sap3/_0103_ heichips25_sap3__3962_/Q
+ heichips25_sap3__4024_/CLK sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm_hold1095 heichips25_can_lehmann_fsm/_0060_ VPWR VGND heichips25_can_lehmann_fsm/net1094
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__2921__652 VPWR VGND net651 sg13g2_tiehi
Xheichips25_sap3__2913_ heichips25_sap3/_0553_ heichips25_sap3/net278 heichips25_sap3/net211
+ VPWR VGND sg13g2_nand2_1
XFILLER_10_985 VPWR VGND sg13g2_decap_8
Xclkload19 VPWR clkload19/Y clkload19/A VGND sg13g2_inv_1
XFILLER_5_455 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3893_ heichips25_sap3/net435 VGND VPWR heichips25_sap3/_0034_ heichips25_sap3__3893_/Q
+ net817 sg13g2_dfrbpq_1
Xheichips25_sap3__2844_ heichips25_sap3/_1869_ heichips25_sap3/_0485_ heichips25_sap3/_0486_
+ heichips25_sap3/_0487_ VPWR VGND sg13g2_nor3_1
XFILLER_5_466 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2775_ heichips25_sap3/_0421_ heichips25_sap3/_0417_ heichips25_sap3/net274
+ heichips25_sap3/_0416_ heichips25_sap3/net288 VPWR VGND sg13g2_a22oi_1
XFILLER_48_153 VPWR VGND sg13g2_decap_4
XFILLER_23_1025 VPWR VGND sg13g2_decap_4
XFILLER_17_540 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3327_ heichips25_sap3/_0937_ heichips25_sap3/net144 heichips25_sap3__3958_/Q
+ heichips25_sap3/net110 heichips25_sap3__3950_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_44_381 VPWR VGND sg13g2_fill_1
XFILLER_44_370 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3258_ heichips25_sap3/_0778_ heichips25_sap3/net53 heichips25_sap3/_0794_
+ heichips25_sap3/_0868_ heichips25_sap3/_0871_ VPWR VGND sg13g2_nor4_1
Xheichips25_sap3__3189_ heichips25_sap3/_0799_ heichips25_sap3/_0800_ heichips25_sap3/_0796_
+ heichips25_sap3/_0802_ VPWR VGND heichips25_sap3/_0801_ sg13g2_nand4_1
Xheichips25_sap3__2209_ heichips25_sap3/_1630_ heichips25_sap3/_1476_ heichips25_sap3/_1496_
+ VPWR VGND sg13g2_nand2_1
XFILLER_20_705 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__3031_ net613 VGND VPWR heichips25_can_lehmann_fsm/net952
+ heichips25_can_lehmann_fsm__3031_/Q clknet_leaf_15_clk sg13g2_dfrbpq_1
XFILLER_39_186 VPWR VGND sg13g2_fill_2
XFILLER_39_164 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2815_ net576 VGND VPWR heichips25_can_lehmann_fsm/_0040_
+ heichips25_can_lehmann_fsm__2815_/Q clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_42_318 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2746_ heichips25_can_lehmann_fsm/net491 VPWR heichips25_can_lehmann_fsm/_0839_
+ VGND heichips25_can_lehmann_fsm/net1127 heichips25_can_lehmann_fsm/net421 sg13g2_o21ai_1
XFILLER_42_329 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2677_ VGND VPWR heichips25_can_lehmann_fsm/_0876_ heichips25_can_lehmann_fsm/net369
+ heichips25_can_lehmann_fsm/_0238_ heichips25_can_lehmann_fsm/_0804_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm_hold915 heichips25_can_lehmann_fsm/_0123_ VPWR VGND heichips25_can_lehmann_fsm/net914
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold904 heichips25_can_lehmann_fsm__2908_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net903 sg13g2_dlygate4sd3_1
XFILLER_10_215 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1628_ VPWR heichips25_can_lehmann_fsm/_0952_ heichips25_can_lehmann_fsm/net1066
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm_hold948 heichips25_can_lehmann_fsm/_0196_ VPWR VGND heichips25_can_lehmann_fsm/net947
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold959 heichips25_can_lehmann_fsm/_0199_ VPWR VGND heichips25_can_lehmann_fsm/net958
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold937 heichips25_can_lehmann_fsm__2930_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net936 sg13g2_dlygate4sd3_1
XFILLER_10_237 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__1559_ VPWR heichips25_can_lehmann_fsm/_0883_ heichips25_can_lehmann_fsm/net844
+ VGND sg13g2_inv_1
XFILLER_2_403 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2875__746 VPWR VGND net745 sg13g2_tiehi
XFILLER_49_11 VPWR VGND sg13g2_decap_8
XFILLER_2_425 VPWR VGND sg13g2_fill_1
XFILLER_2_436 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2560_ heichips25_sap3/_0235_ heichips25_sap3/net77 heichips25_sap3__4022_/Q
+ heichips25_sap3/net90 heichips25_sap3__3942_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2491_ VPWR VGND heichips25_sap3__3972_/Q heichips25_sap3/_1901_
+ heichips25_sap3/net71 heichips25_sap3__4020_/Q heichips25_sap3/_1904_ heichips25_sap3/net79
+ sg13g2_a221oi_1
XFILLER_18_348 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3112_ VGND VPWR heichips25_sap3/_1504_ heichips25_sap3/_1565_ heichips25_sap3/_0725_
+ heichips25_sap3/_1480_ sg13g2_a21oi_1
Xheichips25_sap3__3043_ heichips25_sap3/net238 heichips25_sap3/_1644_ heichips25_sap3/_1449_
+ heichips25_sap3/_0656_ VPWR VGND sg13g2_nand3_1
XFILLER_10_771 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3945_ heichips25_sap3/net444 VGND VPWR heichips25_sap3/_0086_ heichips25_sap3__3945_/Q
+ clkload21/A sg13g2_dfrbpq_1
XFILLER_5_274 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2827_ heichips25_sap3/_0465_ heichips25_sap3/_0466_ heichips25_sap3/_0460_
+ heichips25_sap3/_0471_ VPWR VGND heichips25_sap3/_0470_ sg13g2_nand4_1
Xheichips25_can_lehmann_fsm__2776__655 VPWR VGND net654 sg13g2_tiehi
Xheichips25_sap3__2758_ heichips25_sap3/_0393_ heichips25_sap3/_0377_ heichips25_sap3/_0404_
+ VPWR VGND sg13g2_xor2_1
Xheichips25_sap3__2689_ heichips25_sap3/_1898_ heichips25_sap3/_1877_ heichips25_sap3/_0335_
+ VPWR VGND sg13g2_nor2b_1
XFILLER_49_473 VPWR VGND sg13g2_fill_1
XFILLER_36_101 VPWR VGND sg13g2_fill_1
Xinput6 ui_in[3] net6 VPWR VGND sg13g2_buf_1
XFILLER_36_134 VPWR VGND sg13g2_decap_4
XFILLER_37_679 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2600_ heichips25_can_lehmann_fsm/net493 VPWR heichips25_can_lehmann_fsm/_0766_
+ VGND heichips25_can_lehmann_fsm/net959 heichips25_can_lehmann_fsm/net366 sg13g2_o21ai_1
XFILLER_33_830 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2531_ VGND VPWR heichips25_can_lehmann_fsm/_0915_ heichips25_can_lehmann_fsm/net409
+ heichips25_can_lehmann_fsm/_0165_ heichips25_can_lehmann_fsm/_0731_ sg13g2_a21oi_1
XFILLER_20_524 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2462_ heichips25_can_lehmann_fsm/net499 VPWR heichips25_can_lehmann_fsm/_0697_
+ VGND heichips25_can_lehmann_fsm/net1102 heichips25_can_lehmann_fsm/net429 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2393_ VGND VPWR heichips25_can_lehmann_fsm/_0953_ heichips25_can_lehmann_fsm/net360
+ heichips25_can_lehmann_fsm/_0096_ heichips25_can_lehmann_fsm/_0662_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__3000__594 VPWR VGND net593 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__3014_ net770 VGND VPWR heichips25_can_lehmann_fsm/_0239_
+ heichips25_can_lehmann_fsm__3014_/Q clknet_leaf_19_clk sg13g2_dfrbpq_1
XFILLER_10_38 VPWR VGND sg13g2_fill_2
XFILLER_0_929 VPWR VGND sg13g2_decap_8
XFILLER_16_819 VPWR VGND sg13g2_fill_2
XFILLER_27_145 VPWR VGND sg13g2_decap_8
XFILLER_27_167 VPWR VGND sg13g2_decap_4
XFILLER_42_126 VPWR VGND sg13g2_fill_2
XFILLER_35_35 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2729_ VGND VPWR heichips25_can_lehmann_fsm/_0863_ heichips25_can_lehmann_fsm/net396
+ heichips25_can_lehmann_fsm/_0264_ heichips25_can_lehmann_fsm/_0830_ sg13g2_a21oi_1
XFILLER_23_384 VPWR VGND sg13g2_fill_1
XFILLER_7_528 VPWR VGND sg13g2_decap_8
XFILLER_11_579 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__1991_ VPWR heichips25_sap3/_1417_ heichips25_sap3__3969_/Q VGND
+ sg13g2_inv_1
Xheichips25_sap3__3730_ heichips25_sap3/net1058 heichips25_sap3/_1246_ heichips25_sap3/_1247_
+ VPWR VGND sg13g2_nor2_1
XFILLER_2_200 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__3053__735 VPWR VGND net734 sg13g2_tiehi
Xheichips25_sap3__3661_ VGND VPWR heichips25_sap3/net146 heichips25_sap3/_1206_ heichips25_sap3/_1207_
+ heichips25_sap3/_0889_ sg13g2_a21oi_1
Xheichips25_sap3__3592_ uio_oe_sap3\[6\] net43 heichips25_sap3/_1144_ heichips25_sap3/_1167_
+ VPWR VGND sg13g2_mux2_1
Xheichips25_sap3__2612_ heichips25_sap3/_0283_ heichips25_sap3/_0281_ heichips25_sap3/_0282_
+ heichips25_sap3/_1521_ heichips25_sap3/_1514_ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2543_ heichips25_sap3__3912_/Q heichips25_sap3__3911_/Q heichips25_sap3__3914_/Q
+ heichips25_sap3__3913_/Q heichips25_sap3/_0219_ VPWR VGND sg13g2_nor4_1
XFILLER_47_955 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2474_ heichips25_sap3/_1887_ heichips25_sap3/_1869_ heichips25_sap3/_1886_
+ VPWR VGND sg13g2_nand2_1
XFILLER_18_123 VPWR VGND sg13g2_fill_2
XFILLER_20_1028 VPWR VGND sg13g2_fill_1
XFILLER_34_627 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3026_ VPWR VGND heichips25_sap3/_1541_ heichips25_sap3/_0638_ heichips25_sap3/_1759_
+ heichips25_sap3/_1494_ heichips25_sap3/_0639_ heichips25_sap3/_1626_ sg13g2_a221oi_1
XFILLER_25_90 VPWR VGND sg13g2_fill_1
XFILLER_10_590 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3928_ heichips25_sap3/net436 VGND VPWR heichips25_sap3/_0069_ heichips25_sap3__3928_/Q
+ heichips25_sap3__3988_/CLK sg13g2_dfrbpq_1
Xheichips25_sap3__3859_ VGND VPWR heichips25_sap3/net1071 heichips25_sap3/_1346_ heichips25_sap3/_1356_
+ heichips25_sap3__4047_/Q sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__1962_ heichips25_can_lehmann_fsm/_0323_ heichips25_can_lehmann_fsm/net184
+ heichips25_can_lehmann_fsm/_0321_ heichips25_can_lehmann_fsm/net197 heichips25_can_lehmann_fsm__2779_/Q
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__1893_ VGND VPWR heichips25_can_lehmann_fsm__3049_/Q heichips25_can_lehmann_fsm/_1161_
+ heichips25_can_lehmann_fsm/_1206_ heichips25_can_lehmann_fsm/_1139_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2514_ heichips25_can_lehmann_fsm/net499 VPWR heichips25_can_lehmann_fsm/_0723_
+ VGND heichips25_can_lehmann_fsm/net950 heichips25_can_lehmann_fsm/net426 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2445_ VGND VPWR heichips25_can_lehmann_fsm/_0936_ heichips25_can_lehmann_fsm/net359
+ heichips25_can_lehmann_fsm/_0122_ heichips25_can_lehmann_fsm/_0688_ sg13g2_a21oi_1
XFILLER_21_877 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2376_ heichips25_can_lehmann_fsm/net500 VPWR heichips25_can_lehmann_fsm/_0654_
+ VGND heichips25_can_lehmann_fsm/net983 heichips25_can_lehmann_fsm/net383 sg13g2_o21ai_1
XFILLER_20_376 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_fanout431 heichips25_can_lehmann_fsm/net432 heichips25_can_lehmann_fsm/net431
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout420 heichips25_can_lehmann_fsm/net432 heichips25_can_lehmann_fsm/net420
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout475 heichips25_can_lehmann_fsm/net503 heichips25_can_lehmann_fsm/net475
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout464 heichips25_can_lehmann_fsm/net466 heichips25_can_lehmann_fsm/net464
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout497 heichips25_can_lehmann_fsm/net498 heichips25_can_lehmann_fsm/net497
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout486 heichips25_can_lehmann_fsm/net489 heichips25_can_lehmann_fsm/net486
+ VPWR VGND sg13g2_buf_1
XFILLER_0_759 VPWR VGND sg13g2_fill_1
XFILLER_46_34 VPWR VGND sg13g2_decap_4
XFILLER_46_12 VPWR VGND sg13g2_fill_1
XFILLER_29_977 VPWR VGND sg13g2_decap_4
XFILLER_44_958 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2190_ heichips25_sap3/_1611_ heichips25_sap3/_1596_ heichips25_sap3/_1610_
+ heichips25_sap3/_1594_ heichips25_sap3/_1524_ VPWR VGND sg13g2_a22oi_1
XFILLER_15_104 VPWR VGND sg13g2_decap_8
XFILLER_28_487 VPWR VGND sg13g2_fill_1
XFILLER_44_969 VPWR VGND sg13g2_fill_1
XFILLER_15_137 VPWR VGND sg13g2_decap_8
XFILLER_12_811 VPWR VGND sg13g2_fill_1
XFILLER_31_619 VPWR VGND sg13g2_decap_4
XFILLER_8_804 VPWR VGND sg13g2_decap_4
XFILLER_23_181 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__3020__723 VPWR VGND net722 sg13g2_tiehi
Xheichips25_sap3__1974_ VPWR heichips25_sap3/_1400_ heichips25_sap3__3935_/Q VGND
+ sg13g2_inv_1
Xheichips25_sap3__3713_ uio_oe_sap3\[6\] heichips25_sap3/net114 heichips25_sap3/_1240_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__3644_ heichips25_sap3/_1141_ heichips25_sap3__3993_/Q heichips25_sap3/_1187_
+ heichips25_sap3/_0134_ VPWR VGND sg13g2_mux2_1
Xheichips25_sap3__3575_ heichips25_sap3/net166 heichips25_sap3/_1152_ heichips25_sap3/_1153_
+ heichips25_sap3/_1154_ VPWR VGND sg13g2_nor3_1
XFILLER_23_8 VPWR VGND sg13g2_fill_2
XFILLER_4_1022 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2526_ VGND VPWR heichips25_sap3/net156 heichips25_sap3/_0202_ heichips25_sap3/_0203_
+ heichips25_sap3/_0201_ sg13g2_a21oi_1
XFILLER_35_914 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2457_ heichips25_sap3/net230 heichips25_sap3/_1472_ heichips25_sap3/_1868_
+ heichips25_sap3/_1870_ VPWR VGND sg13g2_a21o_1
XFILLER_19_465 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2388_ heichips25_sap3/_1807_ heichips25_sap3/net80 heichips25_sap3__4025_/Q
+ heichips25_sap3/net84 heichips25_sap3__3961_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__4058_ heichips25_sap3/net453 VGND VPWR heichips25_sap3/_0001_ heichips25_sap3__4058_/Q
+ clknet_leaf_22_clk sg13g2_dfrbpq_1
Xheichips25_sap3__3009_ heichips25_sap3/_0630_ VPWR heichips25_sap3/_0063_ VGND heichips25_sap3/_1399_
+ heichips25_sap3/net202 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2230_ heichips25_can_lehmann_fsm/_1106_ heichips25_can_lehmann_fsm/net1205
+ heichips25_can_lehmann_fsm/_0554_ VPWR VGND sg13g2_xor2_1
Xheichips25_can_lehmann_fsm__2161_ VGND VPWR net11 heichips25_can_lehmann_fsm/_0499_
+ heichips25_can_lehmann_fsm/_0500_ heichips25_can_lehmann_fsm/_0497_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2901__694 VPWR VGND net693 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2092_ heichips25_can_lehmann_fsm/_0433_ heichips25_can_lehmann_fsm/_0432_
+ heichips25_can_lehmann_fsm/net195 heichips25_can_lehmann_fsm/_0434_ VPWR VGND sg13g2_a21o_1
Xheichips25_can_lehmann_fsm__2994_ net641 VGND VPWR heichips25_can_lehmann_fsm/_0219_
+ heichips25_can_lehmann_fsm__2994_/Q clknet_leaf_20_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1945_ VGND VPWR heichips25_can_lehmann_fsm/net1253 heichips25_can_lehmann_fsm/net188
+ heichips25_can_lehmann_fsm/_0308_ heichips25_can_lehmann_fsm/net192 sg13g2_a21oi_1
XFILLER_37_240 VPWR VGND sg13g2_decap_8
XFILLER_26_903 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1876_ heichips25_can_lehmann_fsm/_1190_ heichips25_can_lehmann_fsm/net314
+ heichips25_can_lehmann_fsm__2916_/Q heichips25_can_lehmann_fsm/net318 heichips25_can_lehmann_fsm__2988_/Q
+ VPWR VGND sg13g2_a22oi_1
XFILLER_25_413 VPWR VGND sg13g2_fill_1
XFILLER_21_674 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2428_ heichips25_can_lehmann_fsm/net481 VPWR heichips25_can_lehmann_fsm/_0680_
+ VGND heichips25_can_lehmann_fsm__2888_/Q heichips25_can_lehmann_fsm/net372 sg13g2_o21ai_1
XFILLER_20_162 VPWR VGND sg13g2_fill_1
XFILLER_4_306 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2359_ VGND VPWR heichips25_can_lehmann_fsm/_0962_ heichips25_can_lehmann_fsm/net424
+ heichips25_can_lehmann_fsm/_0079_ heichips25_can_lehmann_fsm/_0645_ sg13g2_a21oi_1
XFILLER_4_317 VPWR VGND sg13g2_fill_1
XFILLER_0_512 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_fanout294 heichips25_can_lehmann_fsm/_1004_ heichips25_can_lehmann_fsm/net294
+ VPWR VGND sg13g2_buf_1
Xheichips25_sap3__3360_ heichips25_sap3/net52 heichips25_sap3/_0922_ heichips25_sap3/net49
+ heichips25_sap3/_0969_ VPWR VGND heichips25_sap3/_0968_ sg13g2_nand4_1
Xheichips25_can_lehmann_fsm__2987__677 VPWR VGND net676 sg13g2_tiehi
Xheichips25_sap3__2311_ heichips25_sap3/_1732_ heichips25_sap3/_1715_ heichips25_sap3/_1730_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__3291_ heichips25_sap3/_0903_ heichips25_sap3/net61 heichips25_sap3/_0852_
+ VPWR VGND sg13g2_xnor2_1
Xheichips25_sap3__2242_ heichips25_sap3/_1507_ VPWR heichips25_sap3/_1663_ VGND heichips25_sap3/_1627_
+ heichips25_sap3/_1662_ sg13g2_o21ai_1
XFILLER_28_251 VPWR VGND sg13g2_decap_4
XFILLER_28_273 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2173_ heichips25_sap3/_1526_ VPWR heichips25_sap3/_1594_ VGND heichips25_sap3/_1499_
+ heichips25_sap3/_1568_ sg13g2_o21ai_1
Xclkbuf_leaf_23_clk clknet_2_0__leaf_clk clknet_leaf_23_clk VPWR VGND sg13g2_buf_8
XFILLER_24_490 VPWR VGND sg13g2_decap_4
Xclkbuf_4_7_0_heichips25_sap3\_sap_3_inst.alu_inst.clk clknet_0_heichips25_sap3\/sap_3_inst.alu_inst.clk
+ clknet_4_7_0_heichips25_sap3\/sap_3_inst.alu_inst.clk VPWR VGND sg13g2_buf_8
XFILLER_7_166 VPWR VGND sg13g2_decap_4
XFILLER_7_155 VPWR VGND sg13g2_fill_2
XFILLER_7_144 VPWR VGND sg13g2_fill_1
XFILLER_7_133 VPWR VGND sg13g2_decap_8
XFILLER_8_689 VPWR VGND sg13g2_decap_8
XFILLER_7_188 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__1957_ VPWR heichips25_sap3/_1383_ heichips25_sap3/net280 VGND sg13g2_inv_1
XFILLER_4_895 VPWR VGND sg13g2_fill_2
XFILLER_4_884 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3627_ heichips25_sap3/_0126_ heichips25_sap3/_1122_ heichips25_sap3/_1185_
+ heichips25_sap3/net103 heichips25_sap3/_1416_ VPWR VGND sg13g2_a22oi_1
XFILLER_39_516 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3558_ heichips25_sap3/_1141_ heichips25_sap3/_1077_ heichips25_sap3/_1079_
+ VPWR VGND sg13g2_nand2b_1
XFILLER_14_4 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2509_ heichips25_sap3/_1908_ heichips25_sap3/_1913_ heichips25_sap3/_1921_
+ uio_out_sap3\[1\] VPWR VGND sg13g2_or3_1
Xheichips25_can_lehmann_fsm__1730_ heichips25_can_lehmann_fsm/_1046_ heichips25_can_lehmann_fsm/_1048_
+ heichips25_can_lehmann_fsm/_0973_ heichips25_can_lehmann_fsm/_1051_ VPWR VGND heichips25_can_lehmann_fsm/_1050_
+ sg13g2_nand4_1
Xheichips25_sap3__3489_ heichips25_sap3/net119 heichips25_sap3/_0860_ heichips25_sap3/_1086_
+ VPWR VGND sg13g2_nor2_1
XFILLER_34_221 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1661_ VPWR heichips25_can_lehmann_fsm/_0985_ net3 VGND
+ sg13g2_inv_1
Xheichips25_can_lehmann_fsm__1592_ VPWR heichips25_can_lehmann_fsm/_0916_ heichips25_can_lehmann_fsm/net1013
+ VGND sg13g2_inv_1
XFILLER_22_449 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_14_clk clknet_2_3__leaf_clk clknet_leaf_14_clk VPWR VGND sg13g2_buf_8
XFILLER_33_1027 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2213_ heichips25_can_lehmann_fsm/_0541_ heichips25_can_lehmann_fsm/net1186
+ heichips25_can_lehmann_fsm/_1103_ VPWR VGND sg13g2_xnor2_1
Xheichips25_can_lehmann_fsm__2144_ heichips25_can_lehmann_fsm/_0483_ heichips25_can_lehmann_fsm/net348
+ heichips25_can_lehmann_fsm__2974_/Q VPWR VGND sg13g2_nand2b_1
Xheichips25_can_lehmann_fsm__2075_ heichips25_can_lehmann_fsm/_0420_ heichips25_can_lehmann_fsm/_0419_
+ heichips25_can_lehmann_fsm/_0418_ VPWR VGND sg13g2_nand2b_1
XFILLER_27_25 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2977_ net716 VGND VPWR heichips25_can_lehmann_fsm/_0202_
+ heichips25_can_lehmann_fsm__2977_/Q clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_26_700 VPWR VGND sg13g2_decap_4
Xheichips25_sap3_fanout132 heichips25_sap3/_0772_ heichips25_sap3/net132 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout121 heichips25_sap3/net122 heichips25_sap3/net121 VPWR VGND
+ sg13g2_buf_1
Xheichips25_can_lehmann_fsm__1928_ heichips25_can_lehmann_fsm/_1237_ heichips25_can_lehmann_fsm/_0289_
+ heichips25_can_lehmann_fsm/_1236_ heichips25_can_lehmann_fsm/_0291_ VPWR VGND heichips25_can_lehmann_fsm/_0290_
+ sg13g2_nand4_1
Xheichips25_sap3_fanout110 heichips25_sap3/_0757_ heichips25_sap3/net110 VPWR VGND
+ sg13g2_buf_1
Xheichips25_can_lehmann_fsm__1859_ net9 heichips25_can_lehmann_fsm/net471 heichips25_can_lehmann_fsm/_1175_
+ VPWR VGND sg13g2_nor2b_1
Xheichips25_sap3_fanout154 heichips25_sap3/_0343_ heichips25_sap3/net154 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout143 heichips25_sap3/_0766_ heichips25_sap3/net143 VPWR VGND
+ sg13g2_buf_1
Xheichips25_can_lehmann_fsm_hold1211 heichips25_can_lehmann_fsm__2807_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1210 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1233 heichips25_can_lehmann_fsm/_0039_ VPWR VGND heichips25_can_lehmann_fsm/net1232
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1200 heichips25_can_lehmann_fsm/_0034_ VPWR VGND heichips25_can_lehmann_fsm/net1199
+ sg13g2_dlygate4sd3_1
XFILLER_43_46 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm_hold1222 heichips25_can_lehmann_fsm__2816_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1221 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1266 heichips25_can_lehmann_fsm/_0024_ VPWR VGND heichips25_can_lehmann_fsm/net1265
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1244 heichips25_can_lehmann_fsm/_0011_ VPWR VGND heichips25_can_lehmann_fsm/net1243
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1255 heichips25_can_lehmann_fsm/_0004_ VPWR VGND heichips25_can_lehmann_fsm/net1254
+ sg13g2_dlygate4sd3_1
Xheichips25_sap3__2860_ VGND VPWR heichips25_sap3/net285 heichips25_sap3/net211 heichips25_sap3/_0502_
+ heichips25_sap3/_0486_ sg13g2_a21oi_1
XFILLER_4_103 VPWR VGND sg13g2_fill_2
XFILLER_4_147 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2791_ heichips25_sap3/_1783_ VPWR heichips25_sap3/_0436_ VGND heichips25_sap3/_1776_
+ heichips25_sap3/_0435_ sg13g2_o21ai_1
XFILLER_49_814 VPWR VGND sg13g2_fill_2
XFILLER_0_353 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3412_ VGND VPWR heichips25_sap3/_0993_ heichips25_sap3/_1015_ heichips25_sap3/_1019_
+ heichips25_sap3/_1018_ sg13g2_a21oi_1
Xheichips25_sap3__3343_ heichips25_sap3/_0943_ VPWR heichips25_sap3/_0953_ VGND heichips25_sap3/_0900_
+ heichips25_sap3/net50 sg13g2_o21ai_1
XFILLER_1_1003 VPWR VGND sg13g2_decap_8
XFILLER_17_722 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2885__726 VPWR VGND net725 sg13g2_tiehi
Xheichips25_sap3__3274_ heichips25_sap3/_0885_ heichips25_sap3/_0886_ heichips25_sap3/_0737_
+ heichips25_sap3/_0887_ VPWR VGND sg13g2_nand3_1
XFILLER_44_552 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2225_ heichips25_sap3/net223 VPWR heichips25_sap3/_1646_ VGND heichips25_sap3/_1619_
+ heichips25_sap3/_1645_ sg13g2_o21ai_1
Xheichips25_sap3__2156_ heichips25_sap3/_1480_ heichips25_sap3/_1516_ heichips25_sap3/_1577_
+ VPWR VGND sg13g2_nor2_1
XFILLER_16_287 VPWR VGND sg13g2_fill_1
XFILLER_31_213 VPWR VGND sg13g2_decap_8
XFILLER_31_257 VPWR VGND sg13g2_fill_1
XFILLER_9_932 VPWR VGND sg13g2_decap_4
XFILLER_12_471 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2087_ heichips25_sap3/_1508_ heichips25_sap3/net261 heichips25_sap3/net262
+ VPWR VGND sg13g2_nand2b_1
Xheichips25_sap3__2989_ heichips25_sap3/_0620_ heichips25_sap3/_0607_ heichips25_sap3__3913_/Q
+ heichips25_sap3/_0606_ heichips25_sap3/_0399_ VPWR VGND sg13g2_a22oi_1
Xclkbuf_leaf_3_clk clknet_2_1__leaf_clk clknet_leaf_3_clk VPWR VGND sg13g2_buf_8
XFILLER_39_313 VPWR VGND sg13g2_fill_2
XFILLER_39_302 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2900_ net695 VGND VPWR heichips25_can_lehmann_fsm/_0125_
+ heichips25_can_lehmann_fsm__2900_/Q clknet_leaf_21_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2831_ net544 VGND VPWR heichips25_can_lehmann_fsm/net1159
+ heichips25_can_lehmann_fsm__2831_/Q clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_47_390 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2762_ heichips25_can_lehmann_fsm/net487 VPWR heichips25_can_lehmann_fsm/_0847_
+ VGND heichips25_can_lehmann_fsm/net1116 heichips25_can_lehmann_fsm/net417 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2786__635 VPWR VGND net634 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__1713_ heichips25_can_lehmann_fsm/_1010_ heichips25_can_lehmann_fsm/_1031_
+ heichips25_can_lehmann_fsm/_1037_ VPWR VGND sg13g2_nor2_1
XFILLER_23_703 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2693_ VGND VPWR heichips25_can_lehmann_fsm/_0872_ heichips25_can_lehmann_fsm/net365
+ heichips25_can_lehmann_fsm/_0246_ heichips25_can_lehmann_fsm/_0812_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__1644_ VPWR heichips25_can_lehmann_fsm/_0968_ heichips25_can_lehmann_fsm/net1088
+ VGND sg13g2_inv_1
XFILLER_35_596 VPWR VGND sg13g2_decap_4
XFILLER_22_213 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__3040__759 VPWR VGND net758 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__1575_ VPWR heichips25_can_lehmann_fsm/_0899_ heichips25_can_lehmann_fsm/net946
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__3003__570 VPWR VGND net569 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2127_ heichips25_can_lehmann_fsm/_0463_ heichips25_can_lehmann_fsm/_0464_
+ heichips25_can_lehmann_fsm/_0462_ heichips25_can_lehmann_fsm/_0466_ VPWR VGND heichips25_can_lehmann_fsm/_0465_
+ sg13g2_nand4_1
XFILLER_1_139 VPWR VGND sg13g2_fill_1
XFILLER_1_117 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2058_ heichips25_can_lehmann_fsm/_0404_ heichips25_can_lehmann_fsm/_0401_
+ heichips25_can_lehmann_fsm/_0405_ heichips25_can_lehmann_fsm/_0406_ VPWR VGND sg13g2_a21o_1
XFILLER_38_35 VPWR VGND sg13g2_decap_4
XFILLER_45_305 VPWR VGND sg13g2_decap_8
XFILLER_45_338 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2010_ VGND VPWR heichips25_sap3/_0018_ heichips25_sap3/_1432_ heichips25_sap3/_1431_
+ sg13g2_or2_1
XFILLER_41_511 VPWR VGND sg13g2_fill_1
XFILLER_13_224 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_hold1041 heichips25_can_lehmann_fsm__2956_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1040 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1030 heichips25_can_lehmann_fsm__3029_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1029 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1052 heichips25_can_lehmann_fsm__3053_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1051 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1063 heichips25_can_lehmann_fsm__2927_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1062 sg13g2_dlygate4sd3_1
Xheichips25_sap3__3961_ heichips25_sap3/net459 VGND VPWR heichips25_sap3/_0102_ heichips25_sap3__3961_/Q
+ heichips25_sap3__3993_/CLK sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm_hold1096 heichips25_can_lehmann_fsm__2881_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1095 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1085 heichips25_can_lehmann_fsm__3054_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1084 sg13g2_dlygate4sd3_1
Xheichips25_sap3__2912_ heichips25_sap3/net211 heichips25_sap3/net281 heichips25_sap3/_0532_
+ heichips25_sap3/_0552_ VPWR VGND sg13g2_a21o_1
XFILLER_5_401 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3892_ heichips25_sap3/net435 VGND VPWR heichips25_sap3/_0033_ heichips25_sap3__3892_/Q
+ net816 sg13g2_dfrbpq_1
Xheichips25_sap3__2843_ heichips25_sap3/_0483_ heichips25_sap3/_0484_ heichips25_sap3/_0486_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__2774_ VGND VPWR heichips25_sap3/net254 heichips25_sap3/net168 heichips25_sap3/_0420_
+ heichips25_sap3/_1888_ sg13g2_a21oi_1
XFILLER_0_161 VPWR VGND sg13g2_fill_1
XFILLER_49_666 VPWR VGND sg13g2_decap_4
XFILLER_49_644 VPWR VGND sg13g2_fill_1
XFILLER_49_677 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3326_ VPWR VGND heichips25_sap3__3998_/Q heichips25_sap3/net128
+ heichips25_sap3/net148 heichips25_sap3__4014_/Q heichips25_sap3/_0936_ heichips25_sap3/net116
+ sg13g2_a221oi_1
Xheichips25_sap3__3257_ heichips25_sap3/net53 heichips25_sap3/_0794_ heichips25_sap3/_0868_
+ heichips25_sap3/_0870_ VPWR VGND sg13g2_nor3_1
Xheichips25_sap3__2208_ heichips25_sap3/_1476_ heichips25_sap3/_1477_ heichips25_sap3/net246
+ heichips25_sap3/_1629_ VPWR VGND sg13g2_nand3_1
Xheichips25_sap3__3188_ heichips25_sap3/_0801_ heichips25_sap3/net144 heichips25_sap3__3968_/Q
+ heichips25_sap3/net129 heichips25_sap3__3944_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_32_566 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2139_ heichips25_sap3/_1560_ heichips25_sap3/_1463_ heichips25_sap3/_1546_
+ VPWR VGND sg13g2_nand2_1
XFILLER_32_577 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__3030_ net629 VGND VPWR heichips25_can_lehmann_fsm/_0255_
+ heichips25_can_lehmann_fsm__3030_/Q clknet_leaf_15_clk sg13g2_dfrbpq_1
XFILLER_28_806 VPWR VGND sg13g2_fill_1
XFILLER_27_316 VPWR VGND sg13g2_fill_2
XFILLER_43_809 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2814_ net578 VGND VPWR heichips25_can_lehmann_fsm/net1232
+ heichips25_can_lehmann_fsm__2814_/Q clknet_leaf_7_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2745_ VGND VPWR heichips25_can_lehmann_fsm/_0859_ heichips25_can_lehmann_fsm/net405
+ heichips25_can_lehmann_fsm/_0272_ heichips25_can_lehmann_fsm/_0838_ sg13g2_a21oi_1
XFILLER_23_511 VPWR VGND sg13g2_fill_1
XFILLER_35_393 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm_hold916 heichips25_can_lehmann_fsm__3010_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net915 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__2676_ heichips25_can_lehmann_fsm/net477 VPWR heichips25_can_lehmann_fsm/_0804_
+ VGND heichips25_can_lehmann_fsm/net923 heichips25_can_lehmann_fsm/net369 sg13g2_o21ai_1
XFILLER_11_706 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_hold905 heichips25_can_lehmann_fsm__2945_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net904 sg13g2_dlygate4sd3_1
XFILLER_23_555 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm_hold949 heichips25_can_lehmann_fsm__2861_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net948 sg13g2_dlygate4sd3_1
XFILLER_10_205 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm_hold938 heichips25_can_lehmann_fsm__2921_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net937 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__1627_ VPWR heichips25_can_lehmann_fsm/_0951_ heichips25_can_lehmann_fsm/net1015
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__1558_ VPWR heichips25_can_lehmann_fsm/_0882_ heichips25_can_lehmann_fsm/net1122
+ VGND sg13g2_inv_1
XFILLER_40_36 VPWR VGND sg13g2_fill_2
XFILLER_49_89 VPWR VGND sg13g2_fill_2
XFILLER_49_67 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2490_ heichips25_sap3/_1903_ heichips25_sap3/net86 heichips25_sap3__3948_/Q
+ heichips25_sap3/net218 heichips25_sap3__4004_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_19_839 VPWR VGND sg13g2_decap_8
XFILLER_46_647 VPWR VGND sg13g2_decap_8
XFILLER_18_327 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3111_ heichips25_sap3/_1565_ heichips25_sap3/_1635_ heichips25_sap3/_0724_
+ VPWR VGND sg13g2_nor2_1
XFILLER_27_872 VPWR VGND sg13g2_decap_4
XFILLER_33_308 VPWR VGND sg13g2_fill_1
XFILLER_41_341 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3042_ heichips25_sap3/_1450_ heichips25_sap3/net234 heichips25_sap3/_1643_
+ heichips25_sap3/_0655_ VPWR VGND sg13g2_nor3_1
Xheichips25_sap3__3944_ heichips25_sap3/net441 VGND VPWR heichips25_sap3/_0085_ heichips25_sap3__3944_/Q
+ heichips25_sap3__4024_/CLK sg13g2_dfrbpq_1
XFILLER_5_231 VPWR VGND sg13g2_fill_2
X_27__513 VPWR VGND net512 sg13g2_tielo
Xheichips25_sap3__2826_ heichips25_sap3/_0470_ heichips25_sap3/_0469_ heichips25_sap3/_0374_
+ heichips25_sap3/_0467_ heichips25_sap3/_0340_ VPWR VGND sg13g2_a22oi_1
XFILLER_2_993 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2757_ heichips25_sap3/_0391_ heichips25_sap3/_0361_ heichips25_sap3/_0403_
+ VPWR VGND sg13g2_xor2_1
Xheichips25_sap3__2688_ heichips25_sap3/_0334_ VPWR heichips25_sap3/_0030_ VGND heichips25_sap3/_1374_
+ heichips25_sap3/net214 sg13g2_o21ai_1
XFILLER_37_625 VPWR VGND sg13g2_decap_4
Xinput7 ui_in[4] net7 VPWR VGND sg13g2_buf_1
Xheichips25_sap3__3309_ heichips25_sap3/_0920_ heichips25_sap3/net105 heichips25_sap3__3941_/Q
+ heichips25_sap3/net108 heichips25_sap3__3949_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_24_308 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2530_ heichips25_can_lehmann_fsm/net478 VPWR heichips25_can_lehmann_fsm/_0731_
+ VGND heichips25_can_lehmann_fsm/net1005 heichips25_can_lehmann_fsm/net410 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2461_ VGND VPWR heichips25_can_lehmann_fsm/_0932_ heichips25_can_lehmann_fsm/net380
+ heichips25_can_lehmann_fsm/_0130_ heichips25_can_lehmann_fsm/_0696_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2392_ heichips25_can_lehmann_fsm/net480 VPWR heichips25_can_lehmann_fsm/_0662_
+ VGND heichips25_can_lehmann_fsm/net1081 heichips25_can_lehmann_fsm/net360 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__3013_ net778 VGND VPWR heichips25_can_lehmann_fsm/_0238_
+ heichips25_can_lehmann_fsm__3013_/Q clknet_leaf_18_clk sg13g2_dfrbpq_1
XFILLER_0_908 VPWR VGND sg13g2_decap_8
XFILLER_19_48 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2911__674 VPWR VGND net673 sg13g2_tiehi
XFILLER_27_124 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2728_ heichips25_can_lehmann_fsm/net465 VPWR heichips25_can_lehmann_fsm/_0830_
+ VGND heichips25_can_lehmann_fsm__3039_/Q heichips25_can_lehmann_fsm/net396 sg13g2_o21ai_1
XFILLER_23_363 VPWR VGND sg13g2_decap_8
XFILLER_24_875 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2659_ VGND VPWR heichips25_can_lehmann_fsm/_0881_ heichips25_can_lehmann_fsm/net428
+ heichips25_can_lehmann_fsm/_0229_ heichips25_can_lehmann_fsm/_0795_ sg13g2_a21oi_1
Xheichips25_sap3__1990_ VPWR heichips25_sap3/_1416_ heichips25_sap3__3985_/Q VGND
+ sg13g2_inv_1
Xheichips25_sap3__3660_ heichips25_sap3/_0943_ heichips25_sap3/_0927_ heichips25_sap3/_1206_
+ VPWR VGND sg13g2_xor2_1
Xheichips25_sap3__2611_ heichips25_sap3/net236 heichips25_sap3/_1584_ heichips25_sap3/_0282_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__3591_ heichips25_sap3/_0109_ heichips25_sap3/_1121_ heichips25_sap3/_1166_
+ heichips25_sap3/net100 heichips25_sap3/_1409_ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2542_ heichips25_sap3__3908_/Q heichips25_sap3__3907_/Q heichips25_sap3__3910_/Q
+ heichips25_sap3__3909_/Q heichips25_sap3/_0218_ VPWR VGND sg13g2_nor4_1
Xheichips25_sap3__2473_ heichips25_sap3/_1880_ heichips25_sap3/_1881_ heichips25_sap3/_1886_
+ VPWR VGND sg13g2_nor2_1
XFILLER_47_934 VPWR VGND sg13g2_fill_1
XFILLER_18_102 VPWR VGND sg13g2_fill_1
XFILLER_19_647 VPWR VGND sg13g2_fill_2
XFILLER_47_989 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2812__583 VPWR VGND net582 sg13g2_tiehi
XFILLER_18_168 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__4074_ heichips25_sap3__4074_/A uo_out_sap3\[5\] VPWR VGND sg13g2_buf_1
Xheichips25_sap3__3025_ VGND VPWR heichips25_sap3/net235 heichips25_sap3/net229 heichips25_sap3/_0638_
+ heichips25_sap3/_1492_ sg13g2_a21oi_1
XFILLER_30_823 VPWR VGND sg13g2_fill_2
XFILLER_14_396 VPWR VGND sg13g2_decap_8
XFILLER_30_856 VPWR VGND sg13g2_fill_2
XFILLER_6_551 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3927_ heichips25_sap3/net436 VGND VPWR heichips25_sap3/_0068_ heichips25_sap3__3927_/Q
+ heichips25_sap3__3927_/CLK sg13g2_dfrbpq_1
XFILLER_6_595 VPWR VGND sg13g2_fill_1
XFILLER_44_4 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3858_ VGND VPWR heichips25_sap3/net342 heichips25_sap3/_1346_ heichips25_sap3/_0187_
+ heichips25_sap3/_1355_ sg13g2_a21oi_1
Xheichips25_sap3__2809_ VPWR VGND heichips25_sap3/_0342_ heichips25_sap3/_0453_ heichips25_sap3/_0448_
+ heichips25_sap3/_0372_ heichips25_sap3/_0454_ heichips25_sap3/_0446_ sg13g2_a221oi_1
Xheichips25_sap3__3789_ heichips25_sap3/_1299_ heichips25_sap3/net293 heichips25_sap3__3989_/Q
+ heichips25_sap3/_1259_ heichips25_sap3__3981_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_38_912 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1961_ VGND VPWR heichips25_can_lehmann_fsm__2781_/Q heichips25_can_lehmann_fsm/net188
+ heichips25_can_lehmann_fsm/_0322_ heichips25_can_lehmann_fsm/net192 sg13g2_a21oi_1
XFILLER_49_282 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1892_ heichips25_can_lehmann_fsm/_1199_ heichips25_can_lehmann_fsm/_1204_
+ heichips25_can_lehmann_fsm/_1162_ heichips25_can_lehmann_fsm/_1205_ VPWR VGND sg13g2_nand3_1
Xheichips25_sap3_hold1106 heichips25_sap3__4055_/Q VPWR VGND heichips25_sap3/net1105
+ sg13g2_dlygate4sd3_1
Xheichips25_sap3_hold1139 heichips25_sap3__4047_/Q VPWR VGND heichips25_sap3/net1138
+ sg13g2_dlygate4sd3_1
XFILLER_21_801 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2513_ VGND VPWR heichips25_can_lehmann_fsm/_0919_ heichips25_can_lehmann_fsm/net386
+ heichips25_can_lehmann_fsm/_0156_ heichips25_can_lehmann_fsm/_0722_ sg13g2_a21oi_1
XFILLER_33_650 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2444_ heichips25_can_lehmann_fsm/net464 VPWR heichips25_can_lehmann_fsm/_0688_
+ VGND heichips25_can_lehmann_fsm/net876 heichips25_can_lehmann_fsm/net357 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2375_ VGND VPWR heichips25_can_lehmann_fsm/_0958_ heichips25_can_lehmann_fsm/net430
+ heichips25_can_lehmann_fsm/_0087_ heichips25_can_lehmann_fsm/_0653_ sg13g2_a21oi_1
XFILLER_21_38 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm_fanout432 heichips25_can_lehmann_fsm/_0623_ heichips25_can_lehmann_fsm/net432
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout421 heichips25_can_lehmann_fsm/net422 heichips25_can_lehmann_fsm/net421
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout410 heichips25_can_lehmann_fsm/net420 heichips25_can_lehmann_fsm/net410
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout465 heichips25_can_lehmann_fsm/net466 heichips25_can_lehmann_fsm/net465
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout498 heichips25_can_lehmann_fsm/net502 heichips25_can_lehmann_fsm/net498
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout476 heichips25_can_lehmann_fsm/net479 heichips25_can_lehmann_fsm/net476
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout487 heichips25_can_lehmann_fsm/net489 heichips25_can_lehmann_fsm/net487
+ VPWR VGND sg13g2_buf_1
XFILLER_47_208 VPWR VGND sg13g2_decap_8
XFILLER_46_79 VPWR VGND sg13g2_fill_2
XFILLER_44_948 VPWR VGND sg13g2_fill_2
XFILLER_44_937 VPWR VGND sg13g2_decap_8
XFILLER_28_477 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2844__808 VPWR VGND net807 sg13g2_tiehi
XFILLER_43_469 VPWR VGND sg13g2_fill_2
XFILLER_11_311 VPWR VGND sg13g2_decap_8
XFILLER_7_315 VPWR VGND sg13g2_decap_8
XFILLER_11_355 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3712_ heichips25_sap3/_0157_ heichips25_sap3/_1121_ heichips25_sap3/_1239_
+ heichips25_sap3/net114 heichips25_sap3/_1405_ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__1973_ VPWR heichips25_sap3/_1399_ heichips25_sap3__3922_/Q VGND
+ sg13g2_inv_1
XFILLER_11_71 VPWR VGND sg13g2_decap_8
XFILLER_11_82 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3643_ VGND VPWR heichips25_sap3/_0869_ heichips25_sap3/_1193_ heichips25_sap3/_1194_
+ heichips25_sap3/_1078_ sg13g2_a21oi_1
XFILLER_39_709 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3574_ uio_oe_sap3\[2\] heichips25_sap3/net95 heichips25_sap3/_1153_
+ VPWR VGND sg13g2_nor2_1
XFILLER_4_1001 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2525_ heichips25_sap3/_0202_ heichips25_sap3__3892_/Q heichips25_sap3/_1788_
+ VPWR VGND sg13g2_nand2_1
XFILLER_35_904 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2456_ VGND VPWR heichips25_sap3/_1472_ heichips25_sap3/net230 heichips25_sap3/_1869_
+ heichips25_sap3/_1868_ sg13g2_a21oi_1
Xheichips25_sap3__2387_ heichips25_sap3/_1806_ heichips25_sap3/net81 heichips25_sap3__3969_/Q
+ heichips25_sap3/net87 heichips25_sap3__3945_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__4057_ heichips25_sap3/net452 VGND VPWR heichips25_sap3/net1020 heichips25_sap3/_0007_
+ clknet_leaf_22_clk sg13g2_dfrbpq_1
XFILLER_15_694 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3008_ heichips25_sap3/_0630_ net47 heichips25_sap3/net202 VPWR VGND
+ sg13g2_nand2_1
XFILLER_14_193 VPWR VGND sg13g2_fill_2
Xinput10 ui_in[7] net10 VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm__2895__706 VPWR VGND net705 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2160_ heichips25_can_lehmann_fsm/_0461_ heichips25_can_lehmann_fsm/net205
+ heichips25_can_lehmann_fsm/_0492_ heichips25_can_lehmann_fsm/_0499_ VPWR VGND sg13g2_nor3_1
Xheichips25_can_lehmann_fsm__2091_ heichips25_can_lehmann_fsm/_0433_ heichips25_can_lehmann_fsm/net199
+ heichips25_can_lehmann_fsm/net1264 heichips25_can_lehmann_fsm/_0304_ heichips25_can_lehmann_fsm/net344
+ VPWR VGND sg13g2_a22oi_1
XFILLER_6_392 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2993_ net649 VGND VPWR heichips25_can_lehmann_fsm/_0218_
+ heichips25_can_lehmann_fsm__2993_/Q clknet_leaf_20_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1944_ heichips25_can_lehmann_fsm/_1235_ heichips25_can_lehmann_fsm/_0303_
+ heichips25_can_lehmann_fsm/_0307_ VPWR VGND sg13g2_nor2_1
Xheichips25_can_lehmann_fsm__1875_ heichips25_can_lehmann_fsm/_1189_ heichips25_can_lehmann_fsm/net307
+ heichips25_can_lehmann_fsm__2940_/Q heichips25_can_lehmann_fsm/net311 heichips25_can_lehmann_fsm__3012_/Q
+ VPWR VGND sg13g2_a22oi_1
XFILLER_26_948 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2427_ VGND VPWR heichips25_can_lehmann_fsm/_0941_ heichips25_can_lehmann_fsm/net413
+ heichips25_can_lehmann_fsm/_0113_ heichips25_can_lehmann_fsm/_0679_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2796__615 VPWR VGND net614 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2358_ heichips25_can_lehmann_fsm/net500 VPWR heichips25_can_lehmann_fsm/_0645_
+ VGND heichips25_can_lehmann_fsm__2854_/Q heichips25_can_lehmann_fsm/net424 sg13g2_o21ai_1
XFILLER_10_1028 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2289_ heichips25_can_lehmann_fsm/net328 VPWR heichips25_can_lehmann_fsm/_0602_
+ VGND heichips25_can_lehmann_fsm/net1209 heichips25_can_lehmann_fsm/net207 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm_fanout295 heichips25_can_lehmann_fsm/_1004_ heichips25_can_lehmann_fsm/net295
+ VPWR VGND sg13g2_buf_1
Xheichips25_sap3__2310_ heichips25_sap3/_1715_ heichips25_sap3/_1730_ heichips25_sap3/_1731_
+ VPWR VGND sg13g2_and2_1
Xheichips25_sap3__3290_ heichips25_sap3/net61 heichips25_sap3/_0852_ heichips25_sap3/_0902_
+ VPWR VGND sg13g2_and2_1
Xheichips25_sap3__2241_ VGND VPWR heichips25_sap3/_1569_ heichips25_sap3/net225 heichips25_sap3/_1662_
+ heichips25_sap3/_1518_ sg13g2_a21oi_1
XFILLER_28_263 VPWR VGND sg13g2_fill_1
XFILLER_29_797 VPWR VGND sg13g2_fill_2
XFILLER_32_907 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2172_ VPWR VGND heichips25_sap3/net247 heichips25_sap3/_1591_ heichips25_sap3/_1566_
+ heichips25_sap3/net249 heichips25_sap3/_1593_ heichips25_sap3/_1469_ sg13g2_a221oi_1
XFILLER_32_918 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2924__640 VPWR VGND net639 sg13g2_tiehi
XFILLER_11_141 VPWR VGND sg13g2_fill_1
XFILLER_40_995 VPWR VGND sg13g2_fill_2
XFILLER_12_697 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__1956_ VPWR heichips25_sap3/_1382_ heichips25_sap3/net278 VGND sg13g2_inv_1
XFILLER_3_373 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3626_ heichips25_sap3/net103 heichips25_sap3/_1078_ heichips25_sap3/_1185_
+ VPWR VGND sg13g2_nor2_1
XFILLER_21_6 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3557_ VGND VPWR heichips25_sap3/net56 heichips25_sap3/_1140_ heichips25_sap3/_0101_
+ heichips25_sap3/_1139_ sg13g2_a21oi_1
Xclkbuf_4_10_0_heichips25_sap3\_sap_3_inst.alu_inst.clk clknet_0_heichips25_sap3\/sap_3_inst.alu_inst.clk
+ clknet_4_10_0_heichips25_sap3\/sap_3_inst.alu_inst.clk VPWR VGND sg13g2_buf_8
Xheichips25_sap3__2508_ VGND VPWR heichips25_sap3/_1916_ heichips25_sap3/_1920_ heichips25_sap3/_1921_
+ heichips25_sap3/net67 sg13g2_a21oi_1
Xheichips25_sap3__3488_ heichips25_sap3/_1085_ heichips25_sap3/net108 heichips25_sap3/_0876_
+ VPWR VGND sg13g2_nand2_1
XFILLER_35_723 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2439_ heichips25_sap3/_1854_ heichips25_sap3__3894_/Q heichips25_sap3/_1788_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_can_lehmann_fsm__1660_ VPWR heichips25_can_lehmann_fsm/_0984_ heichips25_can_lehmann_fsm/net353
+ VGND sg13g2_inv_1
XFILLER_34_255 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1591_ VPWR heichips25_can_lehmann_fsm/_0915_ heichips25_can_lehmann_fsm/net1097
+ VGND sg13g2_inv_1
XFILLER_15_480 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2212_ VGND VPWR heichips25_can_lehmann_fsm/net161 heichips25_can_lehmann_fsm/_0539_
+ heichips25_can_lehmann_fsm/_0037_ heichips25_can_lehmann_fsm/_0540_ sg13g2_a21oi_1
XFILLER_8_72 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2143_ heichips25_can_lehmann_fsm/_0482_ heichips25_can_lehmann_fsm/_0478_
+ heichips25_can_lehmann_fsm/_0481_ heichips25_can_lehmann_fsm/net303 heichips25_can_lehmann_fsm/_0944_
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2074_ heichips25_can_lehmann_fsm/net346 VPWR heichips25_can_lehmann_fsm/_0419_
+ VGND heichips25_can_lehmann_fsm/net1269 heichips25_can_lehmann_fsm/net1274 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2976_ net720 VGND VPWR heichips25_can_lehmann_fsm/net847
+ heichips25_can_lehmann_fsm__2976_/Q clknet_leaf_13_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1927_ heichips25_can_lehmann_fsm/_0290_ heichips25_can_lehmann_fsm/net332
+ heichips25_can_lehmann_fsm__3056_/Q heichips25_can_lehmann_fsm/net297 heichips25_can_lehmann_fsm__2912_/Q
+ VPWR VGND sg13g2_a22oi_1
XFILLER_27_37 VPWR VGND sg13g2_decap_8
Xheichips25_sap3_fanout111 heichips25_sap3/net113 heichips25_sap3/net111 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout100 heichips25_sap3/_0771_ heichips25_sap3/net100 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout122 heichips25_sap3/_0749_ heichips25_sap3/net122 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout144 heichips25_sap3/net145 heichips25_sap3/net144 VPWR VGND
+ sg13g2_buf_1
Xheichips25_can_lehmann_fsm__1858_ VPWR VGND heichips25_can_lehmann_fsm/net1160 heichips25_can_lehmann_fsm/_1173_
+ heichips25_can_lehmann_fsm/_1166_ heichips25_can_lehmann_fsm/_0984_ heichips25_can_lehmann_fsm/_1174_
+ heichips25_can_lehmann_fsm/_1163_ sg13g2_a221oi_1
Xheichips25_sap3_fanout166 heichips25_sap3/_0736_ heichips25_sap3/net166 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout133 heichips25_sap3/_0772_ heichips25_sap3/net133 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout155 heichips25_sap3/net156 heichips25_sap3/net155 VPWR VGND
+ sg13g2_buf_1
Xheichips25_can_lehmann_fsm_hold1212 heichips25_can_lehmann_fsm/_0032_ VPWR VGND heichips25_can_lehmann_fsm/net1211
+ sg13g2_dlygate4sd3_1
XFILLER_43_25 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1789_ heichips25_can_lehmann_fsm/net1217 heichips25_can_lehmann_fsm/net1279
+ heichips25_can_lehmann_fsm/_1104_ heichips25_can_lehmann_fsm/_1105_ VPWR VGND sg13g2_nor3_1
XFILLER_41_759 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm_hold1201 heichips25_can_lehmann_fsm__2830_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1200 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1223 heichips25_can_lehmann_fsm/_0041_ VPWR VGND heichips25_can_lehmann_fsm/net1222
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1267 heichips25_can_lehmann_fsm__2797_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1266 sg13g2_dlygate4sd3_1
XFILLER_43_58 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm_hold1234 heichips25_can_lehmann_fsm__2803_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1233 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1256 heichips25_can_lehmann_fsm__2794_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1255 sg13g2_dlygate4sd3_1
XFILLER_22_962 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_hold1245 heichips25_can_lehmann_fsm__2790_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1244 sg13g2_dlygate4sd3_1
Xheichips25_sap3_hold954 heichips25_sap3__4038_/Q VPWR VGND heichips25_sap3/net953
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1278 heichips25_can_lehmann_fsm__3062_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1277 sg13g2_dlygate4sd3_1
XFILLER_49_1024 VPWR VGND sg13g2_decap_4
XFILLER_4_137 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2790_ heichips25_sap3/_1641_ VPWR heichips25_sap3/_0435_ VGND heichips25_sap3/_1621_
+ heichips25_sap3/_1773_ sg13g2_o21ai_1
XFILLER_0_332 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3411_ heichips25_sap3/net62 heichips25_sap3/_0969_ heichips25_sap3/_1016_
+ heichips25_sap3/_1018_ VPWR VGND sg13g2_nor3_1
Xheichips25_sap3__3342_ heichips25_sap3/_0857_ heichips25_sap3/_0951_ heichips25_sap3/net53
+ heichips25_sap3/_0952_ VPWR VGND sg13g2_nand3_1
XFILLER_16_211 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3273_ heichips25_sap3/_0886_ uio_oe_sap3\[0\] heichips25_sap3/net68
+ VPWR VGND sg13g2_nand2_1
XFILLER_44_564 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2224_ heichips25_sap3/_1645_ heichips25_sap3/net238 heichips25_sap3/_1644_
+ VPWR VGND sg13g2_nand2_1
XFILLER_16_244 VPWR VGND sg13g2_fill_1
XFILLER_16_266 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2155_ VGND VPWR heichips25_sap3/_1458_ heichips25_sap3/_1552_ heichips25_sap3/_1576_
+ heichips25_sap3/_1460_ sg13g2_a21oi_1
XFILLER_16_299 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2086_ heichips25_sap3/net262 heichips25_sap3/net261 heichips25_sap3/_1507_
+ VPWR VGND sg13g2_nor2b_1
XFILLER_8_432 VPWR VGND sg13g2_fill_1
XFILLER_9_966 VPWR VGND sg13g2_fill_2
XFILLER_33_80 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2988_ heichips25_sap3/_0619_ heichips25_sap3/net277 heichips25_sap3/_0605_
+ VPWR VGND sg13g2_nand2_1
XFILLER_3_170 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__1939_ VPWR heichips25_sap3/_1365_ heichips25_sap3/net261 VGND sg13g2_inv_1
Xheichips25_sap3__3609_ heichips25_sap3/_1176_ VPWR heichips25_sap3/_0117_ VGND heichips25_sap3/_1140_
+ heichips25_sap3/net94 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2830_ net546 VGND VPWR heichips25_can_lehmann_fsm/_0055_
+ heichips25_can_lehmann_fsm__2830_/Q clknet_leaf_11_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2761_ VGND VPWR heichips25_can_lehmann_fsm/_0854_ heichips25_can_lehmann_fsm/net376
+ heichips25_can_lehmann_fsm/_0280_ heichips25_can_lehmann_fsm/_0846_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__1712_ VGND VPWR heichips25_can_lehmann_fsm/_1028_ heichips25_can_lehmann_fsm/_1035_
+ heichips25_can_lehmann_fsm/_1036_ heichips25_can_lehmann_fsm/_1022_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2692_ heichips25_can_lehmann_fsm/net473 VPWR heichips25_can_lehmann_fsm/_0812_
+ VGND heichips25_can_lehmann_fsm/net1087 heichips25_can_lehmann_fsm/net364 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__1643_ VPWR heichips25_can_lehmann_fsm/_0967_ heichips25_can_lehmann_fsm/net851
+ VGND sg13g2_inv_1
XFILLER_13_28 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1574_ VPWR heichips25_can_lehmann_fsm/_0898_ heichips25_can_lehmann_fsm/net957
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__2126_ heichips25_can_lehmann_fsm/_0465_ heichips25_can_lehmann_fsm/net295
+ heichips25_can_lehmann_fsm__2976_/Q heichips25_can_lehmann_fsm/net306 heichips25_can_lehmann_fsm__2952_/Q
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2057_ heichips25_can_lehmann_fsm/_0303_ VPWR heichips25_can_lehmann_fsm/_0405_
+ VGND heichips25_can_lehmann_fsm/_0401_ heichips25_can_lehmann_fsm/_0404_ sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2959_ net788 VGND VPWR heichips25_can_lehmann_fsm/_0184_
+ heichips25_can_lehmann_fsm__2959_/Q clknet_leaf_15_clk sg13g2_dfrbpq_1
XFILLER_26_520 VPWR VGND sg13g2_decap_8
XFILLER_14_726 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_hold1031 heichips25_can_lehmann_fsm__2982_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1030 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1075 heichips25_can_lehmann_fsm__3024_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1074 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1042 heichips25_can_lehmann_fsm__2905_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1041 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1064 heichips25_can_lehmann_fsm/_0153_ VPWR VGND heichips25_can_lehmann_fsm/net1063
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1053 heichips25_can_lehmann_fsm/_0278_ VPWR VGND heichips25_can_lehmann_fsm/net1052
+ sg13g2_dlygate4sd3_1
Xheichips25_sap3__3960_ heichips25_sap3/net444 VGND VPWR heichips25_sap3/_0101_ heichips25_sap3__3960_/Q
+ clkload22/A sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm_hold1086 heichips25_can_lehmann_fsm__2863_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1085 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1097 heichips25_can_lehmann_fsm/_0106_ VPWR VGND heichips25_can_lehmann_fsm/net1096
+ sg13g2_dlygate4sd3_1
Xheichips25_sap3__2911_ heichips25_sap3/net65 heichips25_sap3/_0544_ heichips25_sap3/_0550_
+ heichips25_sap3/_0551_ VPWR VGND sg13g2_nor3_1
Xheichips25_sap3__3891_ heichips25_sap3/net447 VGND VPWR heichips25_sap3/_0032_ heichips25_sap3__3891_/Q
+ net815 sg13g2_dfrbpq_1
Xheichips25_sap3__2842_ heichips25_sap3/_0483_ heichips25_sap3/_0484_ heichips25_sap3/_0485_
+ VPWR VGND sg13g2_and2_1
Xheichips25_sap3__2773_ heichips25_sap3/_0419_ heichips25_sap3/net154 heichips25_sap3/_0415_
+ VPWR VGND sg13g2_nand2_1
XFILLER_49_689 VPWR VGND sg13g2_decap_8
XFILLER_17_520 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3325_ heichips25_sap3/_0074_ heichips25_sap3/_0925_ heichips25_sap3/_0932_
+ heichips25_sap3/net55 heichips25_sap3/_1375_ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3256_ heichips25_sap3/_0869_ heichips25_sap3/_0795_ heichips25_sap3/_0868_
+ VPWR VGND sg13g2_nand2b_1
Xheichips25_sap3__2207_ heichips25_sap3/_1441_ heichips25_sap3/_1492_ heichips25_sap3/net244
+ heichips25_sap3/net222 heichips25_sap3/_1628_ VPWR VGND sg13g2_nor4_1
Xheichips25_sap3__3187_ heichips25_sap3/_0800_ heichips25_sap3/net104 heichips25_sap3__3952_/Q
+ heichips25_sap3/net109 heichips25_sap3__3960_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2138_ heichips25_sap3/_1464_ heichips25_sap3/_1547_ heichips25_sap3/_1559_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__2069_ heichips25_sap3/_1490_ heichips25_sap3/net272 heichips25_sap3/net271
+ VPWR VGND sg13g2_nand2b_1
Xheichips25_can_lehmann_fsm__2822__563 VPWR VGND net562 sg13g2_tiehi
XFILLER_5_73 VPWR VGND sg13g2_fill_1
XFILLER_5_95 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2813_ net580 VGND VPWR heichips25_can_lehmann_fsm/net1187
+ heichips25_can_lehmann_fsm__2813_/Q clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_27_339 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2744_ heichips25_can_lehmann_fsm/net474 VPWR heichips25_can_lehmann_fsm/_0838_
+ VGND heichips25_can_lehmann_fsm/net1147 heichips25_can_lehmann_fsm/net405 sg13g2_o21ai_1
XFILLER_35_372 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2675_ VGND VPWR heichips25_can_lehmann_fsm/_0877_ heichips25_can_lehmann_fsm/net416
+ heichips25_can_lehmann_fsm/_0237_ heichips25_can_lehmann_fsm/_0803_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm_hold906 heichips25_can_lehmann_fsm/_0171_ VPWR VGND heichips25_can_lehmann_fsm/net905
+ sg13g2_dlygate4sd3_1
XFILLER_24_38 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm_hold917 heichips25_can_lehmann_fsm__2885_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net916 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold939 heichips25_can_lehmann_fsm/_0146_ VPWR VGND heichips25_can_lehmann_fsm/net938
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold928 heichips25_can_lehmann_fsm__2977_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net927 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__1626_ VPWR heichips25_can_lehmann_fsm/_0950_ heichips25_can_lehmann_fsm/net1110
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__1557_ VPWR heichips25_can_lehmann_fsm/_0881_ heichips25_can_lehmann_fsm/net906
+ VGND sg13g2_inv_1
XFILLER_40_48 VPWR VGND sg13g2_fill_1
XFILLER_2_416 VPWR VGND sg13g2_decap_8
XFILLER_49_46 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2109_ VGND VPWR heichips25_can_lehmann_fsm__3029_/Q heichips25_can_lehmann_fsm/net312
+ heichips25_can_lehmann_fsm/_0448_ heichips25_can_lehmann_fsm/net303 sg13g2_a21oi_1
XFILLER_46_626 VPWR VGND sg13g2_fill_2
XFILLER_18_306 VPWR VGND sg13g2_decap_8
XFILLER_19_818 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3110_ VGND VPWR heichips25_sap3/_1513_ heichips25_sap3/_0722_ heichips25_sap3/_0723_
+ heichips25_sap3/net222 sg13g2_a21oi_1
Xheichips25_sap3__3041_ heichips25_sap3/net234 heichips25_sap3/_1501_ heichips25_sap3/_1506_
+ heichips25_sap3/_0654_ VPWR VGND sg13g2_nor3_1
XFILLER_26_372 VPWR VGND sg13g2_decap_8
XFILLER_14_556 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3943_ heichips25_sap3/net444 VGND VPWR heichips25_sap3/_0084_ heichips25_sap3__3943_/Q
+ heichips25_sap3__4009_/CLK sg13g2_dfrbpq_1
XFILLER_5_221 VPWR VGND sg13g2_fill_1
XFILLER_5_254 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2825_ VGND VPWR heichips25_sap3/_0373_ heichips25_sap3/_0468_ heichips25_sap3/_0469_
+ heichips25_sap3/_0339_ sg13g2_a21oi_1
XFILLER_46_8 VPWR VGND sg13g2_decap_4
XFILLER_2_972 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2756_ VGND VPWR heichips25_sap3/_0402_ heichips25_sap3/_0401_ heichips25_sap3/_0400_
+ sg13g2_or2_1
Xheichips25_sap3__2687_ heichips25_sap3/_0334_ heichips25_sap3__3889_/Q heichips25_sap3/net214
+ VPWR VGND sg13g2_nand2_1
Xinput8 ui_in[5] net8 VPWR VGND sg13g2_buf_1
XFILLER_36_169 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3308_ heichips25_sap3/_0917_ heichips25_sap3/_0918_ heichips25_sap3/_0919_
+ VPWR VGND sg13g2_and2_1
XFILLER_17_361 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3239_ heichips25_sap3/_0850_ heichips25_sap3/_0851_ heichips25_sap3/_0852_
+ VPWR VGND sg13g2_and2_1
XFILLER_32_320 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2460_ heichips25_can_lehmann_fsm/net492 VPWR heichips25_can_lehmann_fsm/_0696_
+ VGND heichips25_can_lehmann_fsm__2904_/Q heichips25_can_lehmann_fsm/net380 sg13g2_o21ai_1
XFILLER_32_364 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2391_ VGND VPWR heichips25_can_lehmann_fsm/_0954_ heichips25_can_lehmann_fsm/net399
+ heichips25_can_lehmann_fsm/_0095_ heichips25_can_lehmann_fsm/_0661_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__3012_ net786 VGND VPWR heichips25_can_lehmann_fsm/_0237_
+ heichips25_can_lehmann_fsm__3012_/Q clknet_leaf_17_clk sg13g2_dfrbpq_1
XFILLER_27_103 VPWR VGND sg13g2_fill_2
XFILLER_28_659 VPWR VGND sg13g2_decap_8
XFILLER_42_106 VPWR VGND sg13g2_fill_1
XFILLER_15_309 VPWR VGND sg13g2_fill_1
XFILLER_35_59 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2727_ VGND VPWR heichips25_can_lehmann_fsm/_0863_ heichips25_can_lehmann_fsm/net361
+ heichips25_can_lehmann_fsm/_0263_ heichips25_can_lehmann_fsm/_0829_ sg13g2_a21oi_1
XFILLER_24_854 VPWR VGND sg13g2_decap_8
XFILLER_23_342 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2658_ heichips25_can_lehmann_fsm/net497 VPWR heichips25_can_lehmann_fsm/_0795_
+ VGND heichips25_can_lehmann_fsm/net920 heichips25_can_lehmann_fsm/net428 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__1609_ VPWR heichips25_can_lehmann_fsm/_0933_ heichips25_can_lehmann_fsm/net996
+ VGND sg13g2_inv_1
XFILLER_11_526 VPWR VGND sg13g2_decap_8
XFILLER_11_537 VPWR VGND sg13g2_fill_1
XFILLER_11_559 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2589_ VGND VPWR heichips25_can_lehmann_fsm/_0900_ heichips25_can_lehmann_fsm/net360
+ heichips25_can_lehmann_fsm/_0194_ heichips25_can_lehmann_fsm/_0760_ sg13g2_a21oi_1
Xheichips25_sap3__2610_ heichips25_sap3/_0281_ heichips25_sap3/_1514_ heichips25_sap3/_1561_
+ VPWR VGND sg13g2_nand2b_1
XFILLER_4_4 VPWR VGND sg13g2_fill_1
XFILLER_2_246 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3590_ heichips25_sap3/_1116_ heichips25_sap3/_1165_ heichips25_sap3/_1166_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__2541_ heichips25_sap3/_0215_ heichips25_sap3/_0216_ heichips25_sap3/_1383_
+ heichips25_sap3/_0217_ VPWR VGND sg13g2_nand3_1
Xheichips25_sap3__2472_ heichips25_sap3/_1880_ heichips25_sap3/_1882_ heichips25_sap3/_1364_
+ heichips25_sap3/_1885_ VPWR VGND sg13g2_nand3_1
Xheichips25_sap3__3872__817 VPWR net816 heichips25_sap3__3927_/CLK VGND sg13g2_inv_1
XFILLER_18_125 VPWR VGND sg13g2_fill_1
XFILLER_20_1019 VPWR VGND sg13g2_decap_8
XFILLER_18_136 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__4073_ heichips25_sap3__4073_/A uo_out_sap3\[4\] VPWR VGND sg13g2_buf_1
XFILLER_33_128 VPWR VGND sg13g2_decap_8
XFILLER_33_139 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3024_ uio_out_sap3\[7\] heichips25_sap3/net259 heichips25_sap3/net231
+ heichips25_sap3/_0071_ VPWR VGND sg13g2_mux2_1
XFILLER_42_695 VPWR VGND sg13g2_fill_1
XFILLER_41_183 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3926_ heichips25_sap3/net436 VGND VPWR heichips25_sap3/_0067_ heichips25_sap3__3926_/Q
+ heichips25_sap3__3927_/CLK sg13g2_dfrbpq_1
Xheichips25_sap3__3857_ heichips25_sap3/net1064 heichips25_sap3/net342 heichips25_sap3/_1355_
+ VPWR VGND sg13g2_nor2_1
XFILLER_37_4 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2808_ heichips25_sap3/_0450_ heichips25_sap3/_0451_ heichips25_sap3/_0447_
+ heichips25_sap3/_0453_ VPWR VGND heichips25_sap3/_0452_ sg13g2_nand4_1
Xheichips25_sap3__3788_ VGND VPWR heichips25_sap3__3941_/Q heichips25_sap3/_1274_
+ heichips25_sap3/_1298_ heichips25_sap3/net290 sg13g2_a21oi_1
XFILLER_2_791 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2739_ heichips25_sap3/net279 heichips25_sap3__3920_/Q heichips25_sap3/_0385_
+ VPWR VGND sg13g2_nor2b_1
Xheichips25_can_lehmann_fsm__1960_ heichips25_can_lehmann_fsm/_0321_ heichips25_can_lehmann_fsm/net1249
+ heichips25_can_lehmann_fsm/_1063_ VPWR VGND sg13g2_xnor2_1
XFILLER_2_30 VPWR VGND sg13g2_fill_2
XFILLER_38_957 VPWR VGND sg13g2_fill_2
XFILLER_2_74 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2969__749 VPWR VGND net748 sg13g2_tiehi
XFILLER_37_467 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1891_ heichips25_can_lehmann_fsm/_1202_ heichips25_can_lehmann_fsm/_1203_
+ heichips25_can_lehmann_fsm/_1201_ heichips25_can_lehmann_fsm/_1204_ VPWR VGND sg13g2_nand3_1
Xheichips25_sap3_hold1129 heichips25_sap3__4032_/Q VPWR VGND heichips25_sap3/net1128
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__2512_ heichips25_can_lehmann_fsm/net499 VPWR heichips25_can_lehmann_fsm/_0722_
+ VGND heichips25_can_lehmann_fsm/net936 heichips25_can_lehmann_fsm/net386 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2443_ VGND VPWR heichips25_can_lehmann_fsm/_0937_ heichips25_can_lehmann_fsm/net394
+ heichips25_can_lehmann_fsm/_0121_ heichips25_can_lehmann_fsm/_0687_ sg13g2_a21oi_1
XFILLER_21_824 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2374_ heichips25_can_lehmann_fsm/net500 VPWR heichips25_can_lehmann_fsm/_0653_
+ VGND heichips25_can_lehmann_fsm/net983 heichips25_can_lehmann_fsm/net430 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm_fanout422 heichips25_can_lehmann_fsm/net425 heichips25_can_lehmann_fsm/net422
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout411 heichips25_can_lehmann_fsm/net420 heichips25_can_lehmann_fsm/net411
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout400 heichips25_can_lehmann_fsm/net408 heichips25_can_lehmann_fsm/net400
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout466 heichips25_can_lehmann_fsm/net470 heichips25_can_lehmann_fsm/net466
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout499 heichips25_can_lehmann_fsm/net502 heichips25_can_lehmann_fsm/net499
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout477 heichips25_can_lehmann_fsm/net478 heichips25_can_lehmann_fsm/net477
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout488 heichips25_can_lehmann_fsm/net489 heichips25_can_lehmann_fsm/net488
+ VPWR VGND sg13g2_buf_1
XFILLER_44_927 VPWR VGND sg13g2_decap_4
XFILLER_11_367 VPWR VGND sg13g2_decap_4
XFILLER_7_349 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3711_ heichips25_sap3/net828 heichips25_sap3/net114 heichips25_sap3/_1116_
+ heichips25_sap3/_1239_ VPWR VGND sg13g2_nor3_1
Xheichips25_sap3__1972_ VPWR heichips25_sap3/_1398_ heichips25_sap3__3921_/Q VGND
+ sg13g2_inv_1
XFILLER_3_544 VPWR VGND sg13g2_decap_4
XFILLER_11_61 VPWR VGND sg13g2_decap_4
XFILLER_11_94 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3642_ VGND VPWR heichips25_sap3/_0794_ heichips25_sap3/_0868_ heichips25_sap3/_1193_
+ heichips25_sap3/_0889_ sg13g2_a21oi_1
Xheichips25_sap3__3573_ net44 heichips25_sap3/net131 heichips25_sap3/_1152_ VPWR VGND
+ sg13g2_nor2_1
Xheichips25_sap3__2524_ heichips25_sap3/net289 heichips25_sap3/net156 heichips25_sap3/_0201_
+ VPWR VGND sg13g2_nor2_1
XFILLER_19_423 VPWR VGND sg13g2_decap_8
XFILLER_46_242 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2455_ heichips25_sap3/_1619_ heichips25_sap3/net221 heichips25_sap3/_1867_
+ heichips25_sap3/_1868_ VPWR VGND sg13g2_nor3_1
XFILLER_47_776 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2386_ heichips25_sap3/_1805_ heichips25_sap3/net72 heichips25_sap3__3977_/Q
+ heichips25_sap3/net216 heichips25_sap3__4009_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_15_640 VPWR VGND sg13g2_fill_2
XFILLER_15_662 VPWR VGND sg13g2_decap_8
XFILLER_15_673 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__4056_ heichips25_sap3/net452 VGND VPWR heichips25_sap3/_0197_ heichips25_sap3__4056_/Q
+ clknet_leaf_23_clk sg13g2_dfrbpq_1
XFILLER_14_150 VPWR VGND sg13g2_fill_2
XFILLER_14_172 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3007_ heichips25_sap3/_0629_ VPWR heichips25_sap3/_0062_ VGND heichips25_sap3/_1398_
+ heichips25_sap3/net202 sg13g2_o21ai_1
Xinput11 uio_in[0] net11 VPWR VGND sg13g2_buf_1
XFILLER_6_360 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2090_ heichips25_can_lehmann_fsm/_0432_ heichips25_can_lehmann_fsm/net186
+ heichips25_can_lehmann_fsm/_0431_ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__3909_ heichips25_sap3/net448 VGND VPWR heichips25_sap3/_0050_ heichips25_sap3__3909_/Q
+ clkload24/A sg13g2_dfrbpq_1
XFILLER_28_0 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2992_ net656 VGND VPWR heichips25_can_lehmann_fsm/_0217_
+ heichips25_can_lehmann_fsm__2992_/Q clknet_leaf_19_clk sg13g2_dfrbpq_1
XFILLER_38_743 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__1943_ VGND VPWR heichips25_can_lehmann_fsm/_1215_ heichips25_can_lehmann_fsm/_0303_
+ heichips25_can_lehmann_fsm/_0306_ heichips25_can_lehmann_fsm/_1234_ sg13g2_a21oi_1
XFILLER_38_798 VPWR VGND sg13g2_fill_1
XFILLER_37_264 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1874_ heichips25_can_lehmann_fsm/_1176_ heichips25_can_lehmann_fsm/_1188_
+ heichips25_can_lehmann_fsm/_0001_ VPWR VGND sg13g2_nor2_1
XFILLER_32_38 VPWR VGND sg13g2_decap_4
XFILLER_20_175 VPWR VGND sg13g2_fill_2
XFILLER_21_687 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2426_ heichips25_can_lehmann_fsm/net481 VPWR heichips25_can_lehmann_fsm/_0679_
+ VGND heichips25_can_lehmann_fsm__2888_/Q heichips25_can_lehmann_fsm/net412 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2357_ VGND VPWR heichips25_can_lehmann_fsm/_0962_ heichips25_can_lehmann_fsm/net383
+ heichips25_can_lehmann_fsm/_0078_ heichips25_can_lehmann_fsm/_0644_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2288_ VGND VPWR heichips25_can_lehmann_fsm/net980 heichips25_can_lehmann_fsm/net171
+ heichips25_can_lehmann_fsm/_0601_ heichips25_can_lehmann_fsm/_0600_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm_fanout296 heichips25_can_lehmann_fsm/net299 heichips25_can_lehmann_fsm/net296
+ VPWR VGND sg13g2_buf_1
XFILLER_29_710 VPWR VGND sg13g2_fill_2
XFILLER_28_220 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2240_ heichips25_sap3/_1661_ heichips25_sap3/_1659_ heichips25_sap3/_1660_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__2171_ heichips25_sap3/_1592_ heichips25_sap3/net247 heichips25_sap3/_1566_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_can_lehmann_fsm__3024__691 VPWR VGND net690 sg13g2_tiehi
XFILLER_7_102 VPWR VGND sg13g2_fill_2
XFILLER_12_676 VPWR VGND sg13g2_decap_4
XFILLER_11_197 VPWR VGND sg13g2_decap_8
XFILLER_22_60 VPWR VGND sg13g2_fill_2
XFILLER_4_831 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__1955_ VPWR heichips25_sap3/_1381_ heichips25_sap3/net286 VGND sg13g2_inv_1
XFILLER_3_341 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3625_ heichips25_sap3/_0125_ heichips25_sap3/_1121_ heichips25_sap3/_1184_
+ heichips25_sap3/net103 heichips25_sap3/_1408_ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3878__823 VPWR net822 heichips25_sap3__3996_/CLK VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__2931__612 VPWR VGND net611 sg13g2_tiehi
Xheichips25_sap3__3556_ heichips25_sap3/_1073_ heichips25_sap3/_1074_ heichips25_sap3/_1140_
+ VPWR VGND sg13g2_nor2_1
XFILLER_14_6 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2507_ heichips25_sap3/_1920_ heichips25_sap3/_1917_ heichips25_sap3/_1918_
+ heichips25_sap3/_1919_ VPWR VGND sg13g2_and3_1
Xheichips25_sap3__3487_ heichips25_sap3/_1084_ heichips25_sap3__3947_/Q heichips25_sap3/net106
+ VPWR VGND sg13g2_nand2_1
XFILLER_19_242 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2438_ VGND VPWR heichips25_sap3/_1853_ heichips25_sap3/net155 heichips25_sap3/net280
+ sg13g2_or2_1
Xheichips25_sap3__2369_ heichips25_sap3/_1790_ heichips25_sap3/net155 heichips25_sap3/_1789_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_can_lehmann_fsm__1590_ VPWR heichips25_can_lehmann_fsm/_0914_ heichips25_can_lehmann_fsm/net970
+ VGND sg13g2_inv_1
XFILLER_34_278 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__4039_ heichips25_sap3/net461 VGND VPWR heichips25_sap3/net1032 heichips25_sap3__4039_/Q
+ clknet_leaf_3_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2211_ heichips25_can_lehmann_fsm/net326 VPWR heichips25_can_lehmann_fsm/_0540_
+ VGND heichips25_can_lehmann_fsm/net1207 heichips25_can_lehmann_fsm/net161 sg13g2_o21ai_1
XFILLER_30_484 VPWR VGND sg13g2_fill_2
XFILLER_30_495 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2142_ VPWR VGND heichips25_can_lehmann_fsm__3052_/Q heichips25_can_lehmann_fsm/_0480_
+ heichips25_can_lehmann_fsm/net333 heichips25_can_lehmann_fsm__2908_/Q heichips25_can_lehmann_fsm/_0481_
+ heichips25_can_lehmann_fsm/net298 sg13g2_a221oi_1
Xheichips25_can_lehmann_fsm__2073_ heichips25_can_lehmann_fsm/net346 heichips25_can_lehmann_fsm/net347
+ heichips25_can_lehmann_fsm/net1274 heichips25_can_lehmann_fsm/_0418_ VPWR VGND sg13g2_nor3_1
XFILLER_6_190 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2832__543 VPWR VGND net542 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2975_ net724 VGND VPWR heichips25_can_lehmann_fsm/_0200_
+ heichips25_can_lehmann_fsm__2975_/Q clknet_leaf_6_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1926_ heichips25_can_lehmann_fsm/_0289_ heichips25_can_lehmann_fsm/net337
+ heichips25_can_lehmann_fsm/_1238_ heichips25_can_lehmann_fsm/net311 heichips25_can_lehmann_fsm__3032_/Q
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3_fanout101 heichips25_sap3/_0771_ heichips25_sap3/net101 VPWR VGND
+ sg13g2_buf_1
XFILLER_38_584 VPWR VGND sg13g2_fill_1
Xheichips25_sap3_fanout123 heichips25_sap3/_0720_ heichips25_sap3/net123 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout112 heichips25_sap3/net113 heichips25_sap3/net112 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout156 heichips25_sap3/_1787_ heichips25_sap3/net156 VPWR VGND
+ sg13g2_buf_1
Xheichips25_can_lehmann_fsm__1857_ heichips25_can_lehmann_fsm/net219 heichips25_can_lehmann_fsm/_1172_
+ heichips25_can_lehmann_fsm/_1173_ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3_fanout134 heichips25_sap3/net137 heichips25_sap3/net134 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout145 heichips25_sap3/_0760_ heichips25_sap3/net145 VPWR VGND
+ sg13g2_buf_1
XFILLER_25_245 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm_hold1213 heichips25_can_lehmann_fsm__2818_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1212 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__1788_ heichips25_can_lehmann_fsm__2813_/Q heichips25_can_lehmann_fsm__2812_/Q
+ heichips25_can_lehmann_fsm__2811_/Q heichips25_can_lehmann_fsm/_1102_ heichips25_can_lehmann_fsm/_1104_
+ VPWR VGND sg13g2_or4_1
Xheichips25_can_lehmann_fsm_hold1202 heichips25_can_lehmann_fsm/_0609_ VPWR VGND heichips25_can_lehmann_fsm/net1201
+ sg13g2_dlygate4sd3_1
Xheichips25_sap3_fanout167 heichips25_sap3/_0605_ heichips25_sap3/net167 VPWR VGND
+ sg13g2_buf_1
X_14__516 VPWR VGND net515 sg13g2_tielo
Xheichips25_can_lehmann_fsm_hold1257 heichips25_can_lehmann_fsm/_0018_ VPWR VGND heichips25_can_lehmann_fsm/net1256
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1246 heichips25_can_lehmann_fsm/_0015_ VPWR VGND heichips25_can_lehmann_fsm/net1245
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1235 heichips25_can_lehmann_fsm__2784_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1234 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1279 heichips25_can_lehmann_fsm__2810_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1278 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1268 heichips25_can_lehmann_fsm/_0023_ VPWR VGND heichips25_can_lehmann_fsm/net1267
+ sg13g2_dlygate4sd3_1
Xheichips25_sap3_hold955 heichips25_sap3/_0179_ VPWR VGND heichips25_sap3/net954 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__2409_ VGND VPWR heichips25_can_lehmann_fsm/_0948_ heichips25_can_lehmann_fsm/net405
+ heichips25_can_lehmann_fsm/_0104_ heichips25_can_lehmann_fsm/_0670_ sg13g2_a21oi_1
XFILLER_49_1003 VPWR VGND sg13g2_decap_8
XFILLER_4_149 VPWR VGND sg13g2_fill_1
XFILLER_4_116 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2993__650 VPWR VGND net649 sg13g2_tiehi
XFILLER_0_311 VPWR VGND sg13g2_fill_1
XFILLER_49_816 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3410_ heichips25_sap3/_0969_ heichips25_sap3/_1016_ heichips25_sap3/_1017_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__3341_ heichips25_sap3/_0777_ heichips25_sap3/net52 heichips25_sap3/net50
+ heichips25_sap3/_0943_ heichips25_sap3/_0951_ VPWR VGND sg13g2_nor4_1
Xheichips25_sap3__3272_ heichips25_sap3/_0885_ uio_out_sap3\[0\] heichips25_sap3/_0884_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__2223_ heichips25_sap3/_1644_ heichips25_sap3/net264 heichips25_sap3/_1441_
+ VPWR VGND sg13g2_nand2_1
XFILLER_44_576 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2154_ VGND VPWR heichips25_sap3/net229 heichips25_sap3/_1553_ heichips25_sap3/_1575_
+ heichips25_sap3/_1513_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2809__589 VPWR VGND net588 sg13g2_tiehi
Xheichips25_sap3__2085_ heichips25_sap3/net258 heichips25_sap3/net260 heichips25_sap3/net267
+ heichips25_sap3/_1506_ VPWR VGND sg13g2_or3_1
XFILLER_9_901 VPWR VGND sg13g2_decap_4
XFILLER_31_248 VPWR VGND sg13g2_decap_8
XFILLER_8_411 VPWR VGND sg13g2_fill_1
XFILLER_12_451 VPWR VGND sg13g2_decap_8
XFILLER_8_444 VPWR VGND sg13g2_decap_8
XFILLER_8_477 VPWR VGND sg13g2_decap_4
XFILLER_8_488 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2987_ VPWR VGND heichips25_sap3/_0408_ heichips25_sap3/_0618_ heichips25_sap3/net153
+ heichips25_sap3/_1382_ heichips25_sap3/_0053_ heichips25_sap3/net167 sg13g2_a221oi_1
Xheichips25_sap3__1938_ VPWR heichips25_sap3/_1364_ heichips25_sap3/net263 VGND sg13g2_inv_1
Xheichips25_sap3__3608_ heichips25_sap3/_1176_ heichips25_sap3__3976_/Q heichips25_sap3/net94
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__3539_ heichips25_sap3/_1129_ heichips25_sap3/net96 heichips25_sap3/_1037_
+ VPWR VGND sg13g2_nand2_1
XFILLER_39_337 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2760_ heichips25_can_lehmann_fsm/net487 VPWR heichips25_can_lehmann_fsm/_0846_
+ VGND heichips25_can_lehmann_fsm__3054_/Q heichips25_can_lehmann_fsm/net376 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__1711_ heichips25_can_lehmann_fsm/_1035_ heichips25_can_lehmann_fsm__3061_/Q
+ heichips25_can_lehmann_fsm/_1034_ VPWR VGND sg13g2_nand2_1
Xheichips25_can_lehmann_fsm__2691_ VGND VPWR heichips25_can_lehmann_fsm/_0873_ heichips25_can_lehmann_fsm/net392
+ heichips25_can_lehmann_fsm/_0245_ heichips25_can_lehmann_fsm/_0811_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__1642_ VPWR heichips25_can_lehmann_fsm/_0966_ heichips25_can_lehmann_fsm/net1006
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__1573_ VPWR heichips25_can_lehmann_fsm/_0897_ heichips25_can_lehmann_fsm/net846
+ VGND sg13g2_inv_1
XFILLER_30_281 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2125_ heichips25_can_lehmann_fsm/_0464_ heichips25_can_lehmann_fsm/net333
+ heichips25_can_lehmann_fsm__3048_/Q heichips25_can_lehmann_fsm/net299 heichips25_can_lehmann_fsm__2904_/Q
+ VPWR VGND sg13g2_a22oi_1
XFILLER_1_119 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2056_ heichips25_can_lehmann_fsm/_0404_ heichips25_can_lehmann_fsm/_0402_
+ heichips25_can_lehmann_fsm/_0403_ VPWR VGND sg13g2_xnor2_1
Xheichips25_can_lehmann_fsm__2958_ net792 VGND VPWR heichips25_can_lehmann_fsm/_0183_
+ heichips25_can_lehmann_fsm__2958_/Q clknet_leaf_15_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1909_ heichips25_can_lehmann_fsm/_1218_ heichips25_can_lehmann_fsm/_1219_
+ heichips25_can_lehmann_fsm/_1217_ heichips25_can_lehmann_fsm/_1222_ VPWR VGND heichips25_can_lehmann_fsm/_1221_
+ sg13g2_nand4_1
Xheichips25_can_lehmann_fsm__2889_ net717 VGND VPWR heichips25_can_lehmann_fsm/net871
+ heichips25_can_lehmann_fsm__2889_/Q clknet_leaf_14_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm_hold1010 heichips25_can_lehmann_fsm/_0126_ VPWR VGND heichips25_can_lehmann_fsm/net1009
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1043 heichips25_can_lehmann_fsm/_0130_ VPWR VGND heichips25_can_lehmann_fsm/net1042
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1054 heichips25_can_lehmann_fsm__2990_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1053 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1087 heichips25_can_lehmann_fsm/_0089_ VPWR VGND heichips25_can_lehmann_fsm/net1086
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1076 heichips25_can_lehmann_fsm/_0250_ VPWR VGND heichips25_can_lehmann_fsm/net1075
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1098 heichips25_can_lehmann_fsm__2939_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1097 sg13g2_dlygate4sd3_1
Xheichips25_sap3__2910_ heichips25_sap3/_0548_ VPWR heichips25_sap3/_0550_ VGND heichips25_sap3/_0341_
+ heichips25_sap3/_0549_ sg13g2_o21ai_1
Xheichips25_sap3__3890_ heichips25_sap3/net447 VGND VPWR heichips25_sap3/_0031_ heichips25_sap3__3890_/Q
+ net814 sg13g2_dfrbpq_1
XFILLER_5_425 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2841_ VGND VPWR heichips25_sap3/net289 heichips25_sap3/_0462_ heichips25_sap3/_0484_
+ heichips25_sap3/_0461_ sg13g2_a21oi_1
Xheichips25_sap3__2772_ heichips25_sap3/_0340_ VPWR heichips25_sap3/_0418_ VGND heichips25_sap3/_0413_
+ heichips25_sap3/_0415_ sg13g2_o21ai_1
XFILLER_49_624 VPWR VGND sg13g2_fill_1
XFILLER_0_174 VPWR VGND sg13g2_decap_4
XFILLER_49_679 VPWR VGND sg13g2_fill_1
XFILLER_37_819 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3324_ heichips25_sap3/_0841_ VPWR heichips25_sap3/_0935_ VGND heichips25_sap3/net61
+ heichips25_sap3/_0852_ sg13g2_o21ai_1
XFILLER_28_70 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3255_ heichips25_sap3/net63 heichips25_sap3/_0820_ heichips25_sap3/_0802_
+ heichips25_sap3/_0868_ VPWR VGND heichips25_sap3/_0864_ sg13g2_nand4_1
Xheichips25_sap3__2206_ heichips25_sap3/_1492_ heichips25_sap3/net222 heichips25_sap3/_1627_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__3186_ heichips25_sap3/_0797_ heichips25_sap3/_0798_ heichips25_sap3/_0799_
+ VPWR VGND sg13g2_and2_1
Xheichips25_sap3__2137_ heichips25_sap3/_1558_ heichips25_sap3/_1530_ heichips25_sap3/net271
+ VPWR VGND sg13g2_nand2b_1
XFILLER_13_760 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2068_ heichips25_sap3/net269 heichips25_sap3/net273 heichips25_sap3/_1489_
+ VPWR VGND sg13g2_nor2b_1
XFILLER_12_292 VPWR VGND sg13g2_decap_8
XFILLER_8_296 VPWR VGND sg13g2_fill_1
Xclkbuf_4_3_0_heichips25_sap3\_sap_3_inst.alu_inst.clk clknet_0_heichips25_sap3\/sap_3_inst.alu_inst.clk
+ clknet_4_3_0_heichips25_sap3\/sap_3_inst.alu_inst.clk VPWR VGND sg13g2_buf_8
XFILLER_39_123 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2812_ net582 VGND VPWR heichips25_can_lehmann_fsm/net1208
+ heichips25_can_lehmann_fsm__2812_/Q clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_27_318 VPWR VGND sg13g2_fill_1
XFILLER_36_852 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2743_ VGND VPWR heichips25_can_lehmann_fsm/_0859_ heichips25_can_lehmann_fsm/net365
+ heichips25_can_lehmann_fsm/_0271_ heichips25_can_lehmann_fsm/_0837_ sg13g2_a21oi_1
XFILLER_36_874 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2674_ heichips25_can_lehmann_fsm/net482 VPWR heichips25_can_lehmann_fsm/_0803_
+ VGND heichips25_can_lehmann_fsm/net923 heichips25_can_lehmann_fsm/net416 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm_hold907 heichips25_can_lehmann_fsm__3003_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net906 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__2983__693 VPWR VGND net692 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__1625_ VPWR heichips25_can_lehmann_fsm/_0949_ heichips25_can_lehmann_fsm/net1126
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm_hold929 heichips25_can_lehmann_fsm__2995_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net928 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold918 heichips25_can_lehmann_fsm/_0111_ VPWR VGND heichips25_can_lehmann_fsm/net917
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__1556_ VPWR heichips25_can_lehmann_fsm/_0880_ heichips25_can_lehmann_fsm/net931
+ VGND sg13g2_inv_1
XFILLER_40_38 VPWR VGND sg13g2_fill_1
XFILLER_49_25 VPWR VGND sg13g2_decap_8
XFILLER_46_1028 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2108_ VGND VPWR heichips25_can_lehmann_fsm/_0445_ heichips25_can_lehmann_fsm/_0446_
+ heichips25_can_lehmann_fsm/_0026_ heichips25_can_lehmann_fsm/_0447_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2039_ heichips25_can_lehmann_fsm/net324 VPWR heichips25_can_lehmann_fsm/_0389_
+ VGND heichips25_can_lehmann_fsm/net1238 heichips25_can_lehmann_fsm/net177 sg13g2_o21ai_1
XFILLER_19_808 VPWR VGND sg13g2_fill_2
XFILLER_27_841 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3040_ heichips25_sap3/_0647_ heichips25_sap3/_0651_ heichips25_sap3/_0643_
+ heichips25_sap3/_0653_ VPWR VGND heichips25_sap3/_0652_ sg13g2_nand4_1
XFILLER_42_855 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2962__777 VPWR VGND net776 sg13g2_tiehi
Xheichips25_sap3__3942_ heichips25_sap3/net456 VGND VPWR heichips25_sap3/_0083_ heichips25_sap3__3942_/Q
+ clkload28/A sg13g2_dfrbpq_1
XFILLER_6_778 VPWR VGND sg13g2_decap_8
XFILLER_5_233 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2824_ heichips25_sap3/_0468_ heichips25_sap3/_0363_ heichips25_sap3/_0364_
+ VPWR VGND sg13g2_xnor2_1
XFILLER_2_951 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2755_ heichips25_sap3/_0401_ heichips25_sap3__3893_/Q heichips25_sap3/_0372_
+ VPWR VGND sg13g2_nand2b_1
XFILLER_7_1000 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2686_ heichips25_sap3/_0333_ VPWR heichips25_sap3/_0029_ VGND heichips25_sap3/_1384_
+ heichips25_sap3/net213 sg13g2_o21ai_1
XFILLER_39_91 VPWR VGND sg13g2_decap_8
XFILLER_49_498 VPWR VGND sg13g2_decap_8
XFILLER_49_487 VPWR VGND sg13g2_fill_1
Xinput9 ui_in[6] net9 VPWR VGND sg13g2_buf_1
XFILLER_36_159 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3307_ heichips25_sap3/_0918_ heichips25_sap3/net137 heichips25_sap3__3965_/Q
+ heichips25_sap3/net138 heichips25_sap3__3973_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3238_ heichips25_sap3/_0842_ heichips25_sap3/_0843_ heichips25_sap3/_0845_
+ heichips25_sap3/_0847_ heichips25_sap3/_0851_ VPWR VGND sg13g2_and4_1
Xheichips25_sap3__3169_ heichips25_sap3/_0780_ heichips25_sap3/_0781_ heichips25_sap3/_0779_
+ heichips25_sap3/_0782_ VPWR VGND sg13g2_nand3_1
Xheichips25_can_lehmann_fsm__2390_ heichips25_can_lehmann_fsm/net480 VPWR heichips25_can_lehmann_fsm/_0661_
+ VGND heichips25_can_lehmann_fsm/net1081 heichips25_can_lehmann_fsm/net399 sg13g2_o21ai_1
XFILLER_9_583 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__3011_ net794 VGND VPWR heichips25_can_lehmann_fsm/net882
+ heichips25_can_lehmann_fsm__3011_/Q clknet_leaf_17_clk sg13g2_dfrbpq_1
XFILLER_42_118 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2726_ heichips25_can_lehmann_fsm/net479 VPWR heichips25_can_lehmann_fsm/_0829_
+ VGND heichips25_can_lehmann_fsm/net848 heichips25_can_lehmann_fsm/net369 sg13g2_o21ai_1
XFILLER_24_833 VPWR VGND sg13g2_decap_8
XFILLER_24_844 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2657_ VGND VPWR heichips25_can_lehmann_fsm/_0881_ heichips25_can_lehmann_fsm/net385
+ heichips25_can_lehmann_fsm/_0228_ heichips25_can_lehmann_fsm/_0794_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2588_ heichips25_can_lehmann_fsm/net476 VPWR heichips25_can_lehmann_fsm/_0760_
+ VGND heichips25_can_lehmann_fsm/net921 heichips25_can_lehmann_fsm/net358 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__1608_ VPWR heichips25_can_lehmann_fsm/_0932_ heichips25_can_lehmann_fsm/net1041
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__1539_ VPWR heichips25_can_lehmann_fsm/_0863_ heichips25_can_lehmann_fsm/net842
+ VGND sg13g2_inv_1
Xheichips25_sap3__2540_ heichips25_sap3/net282 heichips25_sap3/net274 heichips25_sap3/net284
+ heichips25_sap3/net277 heichips25_sap3/_0216_ VPWR VGND sg13g2_nor4_1
XFILLER_47_903 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2471_ heichips25_sap3/_1884_ heichips25_sap3/net263 heichips25_sap3/_1879_
+ VPWR VGND sg13g2_nand2_1
XFILLER_19_616 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__4072_ heichips25_sap3__4072_/A uo_out_sap3\[3\] VPWR VGND sg13g2_buf_1
Xheichips25_sap3__3023_ VGND VPWR heichips25_sap3/_1361_ heichips25_sap3/net231 heichips25_sap3/_0070_
+ heichips25_sap3/_0637_ sg13g2_a21oi_1
XFILLER_6_531 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3925_ heichips25_sap3/net435 VGND VPWR heichips25_sap3/_0066_ heichips25_sap3__3925_/Q
+ heichips25_sap3__3988_/CLK sg13g2_dfrbpq_1
Xheichips25_sap3__3856_ VGND VPWR heichips25_sap3/_1430_ heichips25_sap3/net341 heichips25_sap3/_0186_
+ heichips25_sap3/net830 sg13g2_a21oi_1
XFILLER_44_6 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2807_ heichips25_sap3/_0452_ heichips25_sap3/_0449_ heichips25_sap3/_0364_
+ heichips25_sap3/_0416_ heichips25_sap3/net287 VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3787_ heichips25_sap3/_1297_ heichips25_sap3/_1279_ heichips25_sap3__3965_/Q
+ heichips25_sap3/_1278_ heichips25_sap3__4005_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2738_ heichips25_sap3/_0346_ VPWR heichips25_sap3/_0384_ VGND heichips25_sap3/_0371_
+ heichips25_sap3/_0383_ sg13g2_o21ai_1
XFILLER_49_240 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2669_ VPWR heichips25_sap3/_0328_ uio_oe_sap3\[3\] VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__1890_ VPWR VGND heichips25_can_lehmann_fsm__3055_/Q heichips25_can_lehmann_fsm/_1200_
+ heichips25_can_lehmann_fsm/net332 heichips25_can_lehmann_fsm__3007_/Q heichips25_can_lehmann_fsm/_1203_
+ heichips25_can_lehmann_fsm/net318 sg13g2_a221oi_1
XFILLER_17_170 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2511_ VGND VPWR heichips25_can_lehmann_fsm/_0920_ heichips25_can_lehmann_fsm/net422
+ heichips25_can_lehmann_fsm/_0155_ heichips25_can_lehmann_fsm/_0721_ sg13g2_a21oi_1
XFILLER_33_652 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2442_ heichips25_can_lehmann_fsm/net464 VPWR heichips25_can_lehmann_fsm/_0687_
+ VGND heichips25_can_lehmann_fsm/net876 heichips25_can_lehmann_fsm/net394 sg13g2_o21ai_1
XFILLER_32_173 VPWR VGND sg13g2_fill_2
XFILLER_20_346 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2373_ VGND VPWR heichips25_can_lehmann_fsm/_0958_ heichips25_can_lehmann_fsm/net388
+ heichips25_can_lehmann_fsm/_0086_ heichips25_can_lehmann_fsm/_0652_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm_fanout423 heichips25_can_lehmann_fsm/net425 heichips25_can_lehmann_fsm/net423
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout401 heichips25_can_lehmann_fsm/net402 heichips25_can_lehmann_fsm/net401
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout412 heichips25_can_lehmann_fsm/net414 heichips25_can_lehmann_fsm/net412
+ VPWR VGND sg13g2_buf_1
XFILLER_0_707 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm_fanout478 heichips25_can_lehmann_fsm/net479 heichips25_can_lehmann_fsm/net478
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout467 heichips25_can_lehmann_fsm/net469 heichips25_can_lehmann_fsm/net467
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout489 heichips25_can_lehmann_fsm/net490 heichips25_can_lehmann_fsm/net489
+ VPWR VGND sg13g2_buf_1
XFILLER_28_446 VPWR VGND sg13g2_fill_2
XFILLER_29_969 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2709_ VGND VPWR heichips25_can_lehmann_fsm/_0868_ heichips25_can_lehmann_fsm/net419
+ heichips25_can_lehmann_fsm/_0254_ heichips25_can_lehmann_fsm/_0820_ sg13g2_a21oi_1
XFILLER_23_195 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__1971_ VPWR heichips25_sap3/_1397_ heichips25_sap3__3917_/Q VGND
+ sg13g2_inv_1
Xheichips25_sap3__3710_ heichips25_sap3/_0156_ heichips25_sap3/_1111_ heichips25_sap3/_1238_
+ heichips25_sap3/net114 heichips25_sap3/_1401_ VPWR VGND sg13g2_a22oi_1
XFILLER_3_501 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3641_ heichips25_sap3/_1192_ VPWR heichips25_sap3/_0133_ VGND heichips25_sap3/_1140_
+ heichips25_sap3/_1187_ sg13g2_o21ai_1
XFILLER_3_589 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3572_ heichips25_sap3/_0105_ heichips25_sap3/_1095_ heichips25_sap3/_1151_
+ heichips25_sap3/net100 heichips25_sap3/_1389_ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2523_ net3 heichips25_sap3/_1770_ heichips25_sap3/_0200_ VPWR VGND
+ sg13g2_and2_1
XFILLER_47_766 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2454_ VGND VPWR heichips25_sap3/net238 heichips25_sap3/_1643_ heichips25_sap3/_1867_
+ heichips25_sap3/net227 sg13g2_a21oi_1
Xheichips25_sap3__2385_ heichips25_sap3/_1804_ heichips25_sap3/net73 heichips25_sap3__4001_/Q
+ heichips25_sap3/net77 heichips25_sap3__4017_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__4055_ heichips25_sap3/net451 VGND VPWR heichips25_sap3/_0196_ heichips25_sap3__4055_/Q
+ clknet_leaf_23_clk sg13g2_dfrbpq_1
Xheichips25_sap3__3006_ heichips25_sap3/_0629_ heichips25_sap3/net826 heichips25_sap3/net202
+ VPWR VGND sg13g2_nand2_1
XFILLER_42_493 VPWR VGND sg13g2_fill_1
Xinput12 uio_in[1] net12 VPWR VGND sg13g2_buf_1
XFILLER_30_666 VPWR VGND sg13g2_fill_2
XFILLER_30_699 VPWR VGND sg13g2_decap_4
XFILLER_7_895 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3908_ heichips25_sap3/net447 VGND VPWR heichips25_sap3/_0049_ heichips25_sap3__3908_/Q
+ clkload27/A sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2819__569 VPWR VGND net568 sg13g2_tiehi
Xheichips25_sap3__3839_ heichips25_sap3/_1428_ heichips25_sap3/_0018_ heichips25_sap3/_1343_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_can_lehmann_fsm__2991_ net660 VGND VPWR heichips25_can_lehmann_fsm/net919
+ heichips25_can_lehmann_fsm__2991_/Q clknet_leaf_19_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1942_ heichips25_can_lehmann_fsm/_1215_ heichips25_can_lehmann_fsm/_1235_
+ heichips25_can_lehmann_fsm/_0304_ heichips25_can_lehmann_fsm/_0305_ VPWR VGND sg13g2_nor3_1
XFILLER_37_254 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1873_ heichips25_can_lehmann_fsm/_1187_ VPWR heichips25_can_lehmann_fsm/_1188_
+ VGND heichips25_can_lehmann_fsm/_1165_ heichips25_can_lehmann_fsm/_1186_ sg13g2_o21ai_1
XFILLER_26_939 VPWR VGND sg13g2_fill_2
XFILLER_37_298 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_17_clk clknet_2_2__leaf_clk clknet_leaf_17_clk VPWR VGND sg13g2_buf_8
Xheichips25_can_lehmann_fsm__2843__810 VPWR VGND net809 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2425_ VGND VPWR heichips25_can_lehmann_fsm/_0942_ heichips25_can_lehmann_fsm/net412
+ heichips25_can_lehmann_fsm/_0112_ heichips25_can_lehmann_fsm/_0678_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2356_ heichips25_can_lehmann_fsm/net495 VPWR heichips25_can_lehmann_fsm/_0644_
+ VGND heichips25_can_lehmann_fsm/net911 heichips25_can_lehmann_fsm/net383 sg13g2_o21ai_1
XFILLER_20_198 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2287_ heichips25_can_lehmann_fsm/net171 heichips25_can_lehmann_fsm/_0599_
+ heichips25_can_lehmann_fsm/_0600_ VPWR VGND sg13g2_nor2_1
Xheichips25_can_lehmann_fsm_fanout297 heichips25_can_lehmann_fsm/net299 heichips25_can_lehmann_fsm/net297
+ VPWR VGND sg13g2_buf_1
Xheichips25_sap3__2170_ VGND VPWR heichips25_sap3/_1484_ heichips25_sap3/_1590_ heichips25_sap3/_1591_
+ heichips25_sap3/_1471_ sg13g2_a21oi_1
XFILLER_8_604 VPWR VGND sg13g2_fill_1
XFILLER_22_72 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__1954_ VPWR heichips25_sap3/_1380_ heichips25_sap3__3949_/Q VGND
+ sg13g2_inv_1
XFILLER_4_854 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3624_ heichips25_sap3/net102 heichips25_sap3/_1073_ heichips25_sap3/_1184_
+ VPWR VGND sg13g2_nor2_1
XFILLER_3_397 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3555_ heichips25_sap3__3960_/Q heichips25_sap3/net56 heichips25_sap3/_1139_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__3486_ heichips25_sap3/_1083_ heichips25_sap3__3946_/Q heichips25_sap3/net58
+ heichips25_sap3/_0087_ VPWR VGND sg13g2_mux2_1
Xheichips25_sap3__2506_ heichips25_sap3/_1919_ heichips25_sap3/net82 heichips25_sap3__3972_/Q
+ heichips25_sap3/net86 heichips25_sap3__3956_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_47_552 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2437_ VPWR VGND heichips25_sap3/_1851_ heichips25_sap3/_1654_ heichips25_sap3/_1848_
+ heichips25_sap3/_1400_ heichips25_sap3/_1852_ heichips25_sap3/net90 sg13g2_a221oi_1
XFILLER_35_714 VPWR VGND sg13g2_fill_2
XFILLER_22_408 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2368_ heichips25_sap3/_1789_ heichips25_sap3__3897_/Q heichips25_sap3/_1788_
+ VPWR VGND sg13g2_nand2_1
XFILLER_34_257 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2299_ VGND VPWR heichips25_sap3/_1450_ heichips25_sap3/_1718_ heichips25_sap3/_1720_
+ heichips25_sap3/_1616_ sg13g2_a21oi_1
Xheichips25_sap3__4038_ heichips25_sap3/net460 VGND VPWR heichips25_sap3/net954 heichips25_sap3__4038_/Q
+ clknet_leaf_2_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2210_ heichips25_can_lehmann_fsm/_0539_ heichips25_can_lehmann_fsm/net165
+ heichips25_can_lehmann_fsm/_0538_ heichips25_can_lehmann_fsm/net176 heichips25_can_lehmann_fsm__2844_/Q
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2141_ heichips25_can_lehmann_fsm/_0479_ VPWR heichips25_can_lehmann_fsm/_0480_
+ VGND heichips25_can_lehmann_fsm/_0868_ heichips25_can_lehmann_fsm/_0995_ sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2072_ VPWR VGND heichips25_can_lehmann_fsm/net1266 heichips25_can_lehmann_fsm/net182
+ heichips25_can_lehmann_fsm/net190 heichips25_can_lehmann_fsm/net347 heichips25_can_lehmann_fsm/_0417_
+ heichips25_can_lehmann_fsm/net199 sg13g2_a221oi_1
Xclkbuf_leaf_6_clk clknet_2_1__leaf_clk clknet_leaf_6_clk VPWR VGND sg13g2_buf_8
Xheichips25_can_lehmann_fsm__2974_ net728 VGND VPWR heichips25_can_lehmann_fsm/net958
+ heichips25_can_lehmann_fsm__2974_/Q clknet_leaf_13_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1925_ heichips25_can_lehmann_fsm/_1238_ heichips25_can_lehmann_fsm/net349
+ heichips25_can_lehmann_fsm__2984_/Q VPWR VGND sg13g2_nand2b_1
Xheichips25_sap3_fanout102 heichips25_sap3/_0767_ heichips25_sap3/net102 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout113 heichips25_sap3/_0755_ heichips25_sap3/net113 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout124 heichips25_sap3/net126 heichips25_sap3/net124 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout135 heichips25_sap3/net136 heichips25_sap3/net135 VPWR VGND
+ sg13g2_buf_1
Xheichips25_can_lehmann_fsm__1856_ heichips25_can_lehmann_fsm/_1171_ VPWR heichips25_can_lehmann_fsm/_1172_
+ VGND heichips25_can_lehmann_fsm__2866_/Q heichips25_can_lehmann_fsm/net335 sg13g2_o21ai_1
Xheichips25_sap3_fanout146 heichips25_sap3/net149 heichips25_sap3/net146 VPWR VGND
+ sg13g2_buf_1
Xheichips25_can_lehmann_fsm__1787_ heichips25_can_lehmann_fsm/net1207 heichips25_can_lehmann_fsm__2811_/Q
+ heichips25_can_lehmann_fsm/_1102_ heichips25_can_lehmann_fsm/_1103_ VPWR VGND sg13g2_or3_1
Xheichips25_can_lehmann_fsm_hold1203 heichips25_can_lehmann_fsm__2805_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1202 sg13g2_dlygate4sd3_1
Xheichips25_sap3_fanout168 heichips25_sap3/_1891_ heichips25_sap3/net168 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout157 heichips25_sap3/net158 heichips25_sap3/net157 VPWR VGND
+ sg13g2_buf_1
Xheichips25_can_lehmann_fsm_hold1214 heichips25_can_lehmann_fsm__3063_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1213 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1258 heichips25_can_lehmann_fsm__2782_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1257 sg13g2_dlygate4sd3_1
XFILLER_40_238 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm_hold1236 heichips25_can_lehmann_fsm/_0009_ VPWR VGND heichips25_can_lehmann_fsm/net1235
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1247 heichips25_can_lehmann_fsm__2789_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1246 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1269 heichips25_can_lehmann_fsm__2801_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1268 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__2408_ heichips25_can_lehmann_fsm/net493 VPWR heichips25_can_lehmann_fsm/_0670_
+ VGND heichips25_can_lehmann_fsm/net1000 heichips25_can_lehmann_fsm/net405 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2339_ VGND VPWR heichips25_can_lehmann_fsm/_0967_ heichips25_can_lehmann_fsm/net406
+ heichips25_can_lehmann_fsm/_0069_ heichips25_can_lehmann_fsm/_0635_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2958__793 VPWR VGND net792 sg13g2_tiehi
XFILLER_0_367 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3340_ heichips25_sap3/_0949_ VPWR heichips25_sap3/_0950_ VGND heichips25_sap3/net123
+ heichips25_sap3/_0946_ sg13g2_o21ai_1
Xheichips25_sap3__3271_ heichips25_sap3/_0884_ heichips25_sap3/net127 heichips25_sap3/net131
+ VPWR VGND sg13g2_nand2_1
XFILLER_29_563 VPWR VGND sg13g2_decap_8
XFILLER_44_522 VPWR VGND sg13g2_fill_1
XFILLER_44_511 VPWR VGND sg13g2_decap_8
XFILLER_1_1017 VPWR VGND sg13g2_decap_8
XFILLER_1_1028 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2222_ heichips25_sap3/_1363_ heichips25_sap3/net256 heichips25_sap3/_1643_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__2153_ VPWR heichips25_sap3/_1574_ heichips25_sap3/_1573_ VGND sg13g2_inv_1
Xheichips25_sap3__2084_ heichips25_sap3/net258 heichips25_sap3/net260 heichips25_sap3/net267
+ heichips25_sap3/_1505_ VPWR VGND sg13g2_nor3_1
XFILLER_13_931 VPWR VGND sg13g2_fill_2
XFILLER_31_227 VPWR VGND sg13g2_decap_8
XFILLER_8_423 VPWR VGND sg13g2_decap_8
XFILLER_12_496 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2986_ heichips25_sap3__3912_/Q heichips25_sap3/net167 heichips25_sap3/net153
+ heichips25_sap3/_0618_ VPWR VGND sg13g2_nor3_1
Xheichips25_sap3__1937_ VPWR heichips25_sap3/_1363_ heichips25_sap3/net264 VGND sg13g2_inv_1
XFILLER_3_161 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3607_ heichips25_sap3/_1138_ heichips25_sap3__3975_/Q heichips25_sap3/net94
+ heichips25_sap3/_0116_ VPWR VGND sg13g2_mux2_1
Xheichips25_sap3__3538_ VGND VPWR heichips25_sap3/net54 heichips25_sap3/_0869_ heichips25_sap3/_1128_
+ heichips25_sap3/_1127_ sg13g2_a21oi_1
XFILLER_12_4 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3469_ heichips25_sap3/net98 heichips25_sap3/_0984_ heichips25_sap3/_1069_
+ heichips25_sap3/_1070_ VPWR VGND sg13g2_nor3_1
XFILLER_35_511 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1710_ heichips25_can_lehmann_fsm/_1010_ heichips25_can_lehmann_fsm/_1016_
+ heichips25_can_lehmann_fsm/_1034_ VPWR VGND sg13g2_nor2b_1
Xheichips25_can_lehmann_fsm__2690_ heichips25_can_lehmann_fsm/net469 VPWR heichips25_can_lehmann_fsm/_0811_
+ VGND heichips25_can_lehmann_fsm/net1087 heichips25_can_lehmann_fsm/net392 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__1641_ VPWR heichips25_can_lehmann_fsm/_0965_ heichips25_can_lehmann_fsm/net1050
+ VGND sg13g2_inv_1
XFILLER_35_577 VPWR VGND sg13g2_fill_2
XFILLER_22_205 VPWR VGND sg13g2_fill_2
XFILLER_22_238 VPWR VGND sg13g2_fill_2
XFILLER_22_249 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1572_ VPWR heichips25_can_lehmann_fsm/_0896_ heichips25_can_lehmann_fsm/net927
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__2124_ heichips25_can_lehmann_fsm/_0463_ heichips25_can_lehmann_fsm/net315
+ heichips25_can_lehmann_fsm__2928_/Q heichips25_can_lehmann_fsm/net320 heichips25_can_lehmann_fsm__3000_/Q
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2055_ heichips25_can_lehmann_fsm/_0403_ heichips25_can_lehmann_fsm__2799_/Q
+ heichips25_can_lehmann_fsm/net345 VPWR VGND sg13g2_xnor2_1
XFILLER_38_49 VPWR VGND sg13g2_decap_8
XFILLER_45_319 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2957_ net796 VGND VPWR heichips25_can_lehmann_fsm/net1036
+ heichips25_can_lehmann_fsm__2957_/Q clknet_leaf_15_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1908_ heichips25_can_lehmann_fsm/_1221_ heichips25_can_lehmann_fsm/_1220_
+ heichips25_can_lehmann_fsm/net337 heichips25_can_lehmann_fsm/net297 heichips25_can_lehmann_fsm__2913_/Q
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2888_ net719 VGND VPWR heichips25_can_lehmann_fsm/net1004
+ heichips25_can_lehmann_fsm__2888_/Q clknet_leaf_14_clk sg13g2_dfrbpq_1
XFILLER_26_555 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1839_ heichips25_can_lehmann_fsm/_1155_ heichips25_can_lehmann_fsm/net348
+ heichips25_can_lehmann_fsm__3060_/Q VPWR VGND sg13g2_nand2b_1
Xheichips25_can_lehmann_fsm_hold1022 heichips25_can_lehmann_fsm__2989_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1021 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1000 heichips25_can_lehmann_fsm/_0242_ VPWR VGND heichips25_can_lehmann_fsm/net999
+ sg13g2_dlygate4sd3_1
XFILLER_13_249 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm_hold1011 heichips25_can_lehmann_fsm__2994_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1010 sg13g2_dlygate4sd3_1
XFILLER_10_901 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm_hold1044 heichips25_can_lehmann_fsm__3055_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1043 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1055 heichips25_can_lehmann_fsm__2924_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1054 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1077 heichips25_can_lehmann_fsm__3025_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1076 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1099 heichips25_can_lehmann_fsm/_0164_ VPWR VGND heichips25_can_lehmann_fsm/net1098
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1088 heichips25_can_lehmann_fsm__3020_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1087 sg13g2_dlygate4sd3_1
XFILLER_10_967 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2840_ heichips25_sap3/_0483_ heichips25_sap3/net285 heichips25_sap3/net212
+ VPWR VGND sg13g2_xnor2_1
XFILLER_5_448 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2771_ heichips25_sap3/net169 heichips25_sap3/_1896_ heichips25_sap3/_0417_
+ VPWR VGND sg13g2_nor2b_1
XFILLER_0_142 VPWR VGND sg13g2_decap_4
XFILLER_48_157 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3323_ heichips25_sap3/net61 heichips25_sap3/_0865_ heichips25_sap3/_0934_
+ VPWR VGND sg13g2_nor2_1
XFILLER_28_60 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3254_ heichips25_sap3/_0820_ heichips25_sap3/_0864_ heichips25_sap3/net63
+ heichips25_sap3/_0867_ VPWR VGND sg13g2_nand3_1
XFILLER_17_555 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3185_ heichips25_sap3/_0798_ heichips25_sap3/net135 heichips25_sap3__3976_/Q
+ heichips25_sap3/net142 heichips25_sap3__3992_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2205_ VPWR heichips25_sap3/_1626_ heichips25_sap3/net222 VGND sg13g2_inv_1
Xheichips25_sap3__2136_ heichips25_sap3/net267 heichips25_sap3/net269 heichips25_sap3/_1529_
+ heichips25_sap3/_1557_ VPWR VGND sg13g2_nor3_1
Xheichips25_sap3__2067_ heichips25_sap3/_1488_ heichips25_sap3/net258 heichips25_sap3/net260
+ VPWR VGND sg13g2_nand2_1
XFILLER_12_260 VPWR VGND sg13g2_fill_1
XFILLER_8_286 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2969_ heichips25_sap3/_1883_ heichips25_sap3/_1893_ heichips25_sap3/_0606_
+ VPWR VGND sg13g2_nor2_1
XFILLER_4_492 VPWR VGND sg13g2_fill_2
XFILLER_39_102 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2811_ net584 VGND VPWR heichips25_can_lehmann_fsm/_0036_
+ heichips25_can_lehmann_fsm__2811_/Q clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_39_157 VPWR VGND sg13g2_decap_8
XFILLER_39_135 VPWR VGND sg13g2_fill_2
XFILLER_39_179 VPWR VGND sg13g2_decap_8
XFILLER_35_341 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2742_ heichips25_can_lehmann_fsm/net472 VPWR heichips25_can_lehmann_fsm/_0837_
+ VGND heichips25_can_lehmann_fsm/net1154 heichips25_can_lehmann_fsm/net365 sg13g2_o21ai_1
XFILLER_36_886 VPWR VGND sg13g2_fill_2
XFILLER_35_363 VPWR VGND sg13g2_decap_4
XFILLER_35_352 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2673_ VGND VPWR heichips25_can_lehmann_fsm/_0877_ heichips25_can_lehmann_fsm/net374
+ heichips25_can_lehmann_fsm/_0236_ heichips25_can_lehmann_fsm/_0802_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm_hold908 heichips25_can_lehmann_fsm/_0228_ VPWR VGND heichips25_can_lehmann_fsm/net907
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__1624_ VPWR heichips25_can_lehmann_fsm/_0948_ heichips25_can_lehmann_fsm/net1055
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm_hold919 heichips25_can_lehmann_fsm__2991_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net918 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__3044__695 VPWR VGND net694 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__1555_ VPWR heichips25_can_lehmann_fsm/_0879_ heichips25_can_lehmann_fsm/net1139
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__2801__605 VPWR VGND net604 sg13g2_tiehi
XFILLER_31_591 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2107_ heichips25_can_lehmann_fsm/net323 VPWR heichips25_can_lehmann_fsm/_0447_
+ VGND heichips25_can_lehmann_fsm/net1268 heichips25_can_lehmann_fsm/net180 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2990__665 VPWR VGND net664 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2038_ heichips25_can_lehmann_fsm/_0387_ heichips25_can_lehmann_fsm/_0385_
+ heichips25_can_lehmann_fsm/_0386_ heichips25_can_lehmann_fsm/_0388_ VPWR VGND sg13g2_a21o_1
Xheichips25_can_lehmann_fsm__2851__794 VPWR VGND net793 sg13g2_tiehi
XFILLER_41_311 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__3062__751 VPWR VGND net750 sg13g2_tiehi
XFILLER_41_355 VPWR VGND sg13g2_decap_8
XFILLER_41_399 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3941_ heichips25_sap3/net456 VGND VPWR heichips25_sap3/_0082_ heichips25_sap3__3941_/Q
+ heichips25_sap3__4021_/CLK sg13g2_dfrbpq_1
XFILLER_10_786 VPWR VGND sg13g2_fill_2
XFILLER_5_267 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2823_ heichips25_sap3/_0467_ heichips25_sap3/_0400_ heichips25_sap3/_0401_
+ VPWR VGND sg13g2_xnor2_1
XFILLER_30_72 VPWR VGND sg13g2_decap_8
XFILLER_2_930 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2754_ heichips25_sap3/_0389_ heichips25_sap3/_0363_ heichips25_sap3/_0400_
+ VPWR VGND sg13g2_xor2_1
Xheichips25_sap3__2685_ heichips25_sap3/_0333_ heichips25_sap3__3888_/Q heichips25_sap3/net213
+ VPWR VGND sg13g2_nand2_1
XFILLER_36_138 VPWR VGND sg13g2_fill_2
XFILLER_18_831 VPWR VGND sg13g2_fill_2
XFILLER_18_842 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3306_ heichips25_sap3/_0917_ heichips25_sap3/net133 heichips25_sap3__3989_/Q
+ heichips25_sap3/net140 heichips25_sap3__3981_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_18_875 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3237_ heichips25_sap3/_0844_ heichips25_sap3/_0846_ heichips25_sap3/_0848_
+ heichips25_sap3/_0849_ heichips25_sap3/_0850_ VPWR VGND sg13g2_and4_1
Xheichips25_sap3__3168_ heichips25_sap3/_0781_ heichips25_sap3/net132 heichips25_sap3__4002_/Q
+ heichips25_sap3/net142 heichips25_sap3__3994_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2119_ heichips25_sap3/_1540_ heichips25_sap3/_1538_ heichips25_sap3/_1500_
+ VPWR VGND sg13g2_nand2b_1
Xheichips25_sap3__3099_ VPWR VGND heichips25_sap3/_1526_ heichips25_sap3/_0710_ heichips25_sap3/_0711_
+ heichips25_sap3/_1524_ heichips25_sap3/_0712_ heichips25_sap3/_1534_ sg13g2_a221oi_1
Xheichips25_can_lehmann_fsm__3010_ net802 VGND VPWR heichips25_can_lehmann_fsm/_0235_
+ heichips25_can_lehmann_fsm__3010_/Q clknet_leaf_17_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__3039__775 VPWR VGND net774 sg13g2_tiehi
XFILLER_27_105 VPWR VGND sg13g2_fill_1
XFILLER_27_138 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2725_ VGND VPWR heichips25_can_lehmann_fsm/_0864_ heichips25_can_lehmann_fsm/net410
+ heichips25_can_lehmann_fsm/_0262_ heichips25_can_lehmann_fsm/_0828_ sg13g2_a21oi_1
XFILLER_24_812 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2829__549 VPWR VGND net548 sg13g2_tiehi
XFILLER_23_344 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2656_ heichips25_can_lehmann_fsm/net497 VPWR heichips25_can_lehmann_fsm/_0794_
+ VGND heichips25_can_lehmann_fsm__3002_/Q heichips25_can_lehmann_fsm/net385 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2587_ VGND VPWR heichips25_can_lehmann_fsm/_0901_ heichips25_can_lehmann_fsm/net396
+ heichips25_can_lehmann_fsm/_0193_ heichips25_can_lehmann_fsm/_0759_ sg13g2_a21oi_1
XFILLER_23_377 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1607_ VPWR heichips25_can_lehmann_fsm/_0931_ heichips25_can_lehmann_fsm/net900
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__1538_ VPWR heichips25_can_lehmann_fsm/_0862_ heichips25_can_lehmann_fsm/net944
+ VGND sg13g2_inv_1
XFILLER_2_226 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2470_ heichips25_sap3/_1883_ heichips25_sap3/_1880_ heichips25_sap3/_1882_
+ VPWR VGND sg13g2_nand2_1
XFILLER_19_606 VPWR VGND sg13g2_decap_4
XFILLER_18_116 VPWR VGND sg13g2_decap_8
XFILLER_47_959 VPWR VGND sg13g2_fill_1
XFILLER_42_631 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__4071_ heichips25_sap3__4071_/A uo_out_sap3\[2\] VPWR VGND sg13g2_buf_1
Xheichips25_sap3__3022_ heichips25_sap3/net231 heichips25_sap3/net826 heichips25_sap3/_0637_
+ VPWR VGND sg13g2_nor2_1
XFILLER_15_867 VPWR VGND sg13g2_decap_4
XFILLER_41_152 VPWR VGND sg13g2_fill_2
XFILLER_6_510 VPWR VGND sg13g2_decap_8
XFILLER_10_572 VPWR VGND sg13g2_decap_4
XFILLER_41_82 VPWR VGND sg13g2_fill_2
XFILLER_41_60 VPWR VGND sg13g2_fill_1
XFILLER_6_543 VPWR VGND sg13g2_fill_2
XFILLER_10_594 VPWR VGND sg13g2_fill_1
XFILLER_10_583 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3924_ heichips25_sap3/net435 VGND VPWR heichips25_sap3/_0065_ heichips25_sap3__3924_/Q
+ heichips25_sap3__4005_/CLK sg13g2_dfrbpq_1
Xheichips25_sap3__3855_ VGND VPWR heichips25_sap3/_1346_ heichips25_sap3/_1354_ heichips25_sap3/_0185_
+ heichips25_sap3/_1347_ sg13g2_a21oi_1
Xheichips25_sap3__2806_ heichips25_sap3/_1894_ heichips25_sap3/_1896_ heichips25_sap3/net254
+ heichips25_sap3/_0451_ VPWR VGND sg13g2_nand3_1
Xheichips25_can_lehmann_fsm__2934__600 VPWR VGND net599 sg13g2_tiehi
Xheichips25_sap3__3786_ heichips25_sap3/_1296_ heichips25_sap3/_1282_ heichips25_sap3__3949_/Q
+ heichips25_sap3/net292 heichips25_sap3__3957_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_37_6 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2737_ heichips25_sap3/_0355_ heichips25_sap3/_0379_ heichips25_sap3/_0382_
+ heichips25_sap3/_0383_ VPWR VGND sg13g2_nor3_1
Xheichips25_sap3__2668_ VPWR VGND heichips25_sap3/_0231_ heichips25_sap3/net66 heichips25_sap3/_0227_
+ heichips25_sap3/_1368_ uio_oe_sap3\[3\] heichips25_sap3/net92 sg13g2_a221oi_1
XFILLER_49_252 VPWR VGND sg13g2_decap_8
XFILLER_49_296 VPWR VGND sg13g2_decap_8
XFILLER_38_959 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2599_ heichips25_sap3/net280 heichips25_sap3/net279 heichips25_sap3/_0271_
+ VPWR VGND sg13g2_xor2_1
Xheichips25_can_lehmann_fsm__2510_ heichips25_can_lehmann_fsm/net499 VPWR heichips25_can_lehmann_fsm/_0721_
+ VGND heichips25_can_lehmann_fsm/net936 heichips25_can_lehmann_fsm/net422 sg13g2_o21ai_1
XFILLER_36_1028 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2441_ VGND VPWR heichips25_can_lehmann_fsm/_0937_ heichips25_can_lehmann_fsm/net357
+ heichips25_can_lehmann_fsm/_0120_ heichips25_can_lehmann_fsm/_0686_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2372_ heichips25_can_lehmann_fsm/net501 VPWR heichips25_can_lehmann_fsm/_0652_
+ VGND heichips25_can_lehmann_fsm__2860_/Q heichips25_can_lehmann_fsm/net388 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm_fanout424 heichips25_can_lehmann_fsm/net425 heichips25_can_lehmann_fsm/net424
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout402 heichips25_can_lehmann_fsm/net403 heichips25_can_lehmann_fsm/net402
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout413 heichips25_can_lehmann_fsm/net414 heichips25_can_lehmann_fsm/net413
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout479 heichips25_can_lehmann_fsm/net490 heichips25_can_lehmann_fsm/net479
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout468 heichips25_can_lehmann_fsm/net469 heichips25_can_lehmann_fsm/net468
+ VPWR VGND sg13g2_buf_1
XFILLER_46_49 VPWR VGND sg13g2_fill_1
XFILLER_46_38 VPWR VGND sg13g2_fill_1
XFILLER_37_970 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__3007__538 VPWR VGND net537 sg13g2_tiehi
XFILLER_12_804 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2708_ heichips25_can_lehmann_fsm/net486 VPWR heichips25_can_lehmann_fsm/_0820_
+ VGND heichips25_can_lehmann_fsm/net1029 heichips25_can_lehmann_fsm/net419 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2639_ VGND VPWR heichips25_can_lehmann_fsm/_0888_ heichips25_can_lehmann_fsm/net398
+ heichips25_can_lehmann_fsm/_0219_ heichips25_can_lehmann_fsm/_0785_ sg13g2_a21oi_1
XFILLER_8_808 VPWR VGND sg13g2_fill_1
XFILLER_7_329 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__1970_ VPWR heichips25_sap3/_1396_ heichips25_sap3__3916_/Q VGND
+ sg13g2_inv_1
XFILLER_11_41 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3640_ heichips25_sap3/_1192_ heichips25_sap3__3992_/Q heichips25_sap3/net93
+ VPWR VGND sg13g2_nand2_1
XFILLER_3_557 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3571_ heichips25_sap3/net100 heichips25_sap3/_1150_ heichips25_sap3/_1151_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__2522_ VPWR VGND heichips25_sap3/_0198_ heichips25_sap3/_1654_ heichips25_sap3/_1930_
+ heichips25_sap3/_1392_ heichips25_sap3/_0199_ heichips25_sap3/net89 sg13g2_a221oi_1
Xheichips25_sap3__2453_ heichips25_sap3/_1865_ heichips25_sap3/net224 heichips25_sap3/net221
+ heichips25_sap3/_1866_ VPWR VGND sg13g2_a21o_1
XFILLER_4_1015 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2384_ heichips25_sap3__3937_/Q heichips25_sap3/_1734_ heichips25_sap3/_1803_
+ VPWR VGND sg13g2_nor2_1
XFILLER_19_469 VPWR VGND sg13g2_fill_1
XFILLER_28_981 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__4054_ heichips25_sap3/net452 VGND VPWR heichips25_sap3/net1125 heichips25_sap3__4054_/Q
+ clknet_leaf_23_clk sg13g2_dfrbpq_1
XFILLER_15_642 VPWR VGND sg13g2_fill_1
XFILLER_14_152 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3005_ heichips25_sap3__3920_/Q uio_out_sap3\[5\] heichips25_sap3/net202
+ heichips25_sap3/_0061_ VPWR VGND sg13g2_mux2_1
XFILLER_30_645 VPWR VGND sg13g2_decap_4
Xinput13 uio_in[2] net13 VPWR VGND sg13g2_buf_1
XFILLER_7_852 VPWR VGND sg13g2_fill_2
XFILLER_7_841 VPWR VGND sg13g2_fill_2
XFILLER_10_380 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3907_ heichips25_sap3/net447 VGND VPWR heichips25_sap3/_0048_ heichips25_sap3__3907_/Q
+ heichips25_sap3__3927_/CLK sg13g2_dfrbpq_1
Xheichips25_sap3__3838_ heichips25_sap3/_0008_ heichips25_sap3/net1031 heichips25_sap3/_1342_
+ heichips25_sap3/_0180_ VPWR VGND sg13g2_a21o_1
Xheichips25_sap3__3769_ heichips25_sap3/_1258_ heichips25_sap3/_1264_ heichips25_sap3/_1281_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3_sap_3_inst.clock.clock_gate_inst heichips25_sap3/_0002_ heichips25_sap3/clk_div_out
+ heichips25_sap3/sap_3_inst.alu_inst.clk VPWR VGND sg13g2_lgcp_1
Xheichips25_can_lehmann_fsm__2990_ net664 VGND VPWR heichips25_can_lehmann_fsm/_0215_
+ heichips25_can_lehmann_fsm__2990_/Q clknet_leaf_19_clk sg13g2_dfrbpq_1
XFILLER_28_2 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1941_ heichips25_can_lehmann_fsm/_0294_ heichips25_can_lehmann_fsm/_0293_
+ heichips25_can_lehmann_fsm/_0302_ heichips25_can_lehmann_fsm/_0304_ VPWR VGND sg13g2_a21o_1
Xheichips25_can_lehmann_fsm__1872_ heichips25_can_lehmann_fsm/_1187_ heichips25_can_lehmann_fsm/_1165_
+ heichips25_can_lehmann_fsm/net352 VPWR VGND sg13g2_nand2b_1
XFILLER_25_406 VPWR VGND sg13g2_decap_8
Xheichips25_sap3_fanout339 heichips25_sap3/net340 heichips25_sap3/net339 VPWR VGND
+ sg13g2_buf_1
XFILLER_20_133 VPWR VGND sg13g2_fill_2
XFILLER_21_667 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2424_ heichips25_can_lehmann_fsm/net481 VPWR heichips25_can_lehmann_fsm/_0678_
+ VGND heichips25_can_lehmann_fsm/net1003 heichips25_can_lehmann_fsm/net412 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2355_ VGND VPWR heichips25_can_lehmann_fsm/_0963_ heichips25_can_lehmann_fsm/net423
+ heichips25_can_lehmann_fsm/_0077_ heichips25_can_lehmann_fsm/_0643_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm_fanout210 heichips25_can_lehmann_fsm/_0476_ heichips25_can_lehmann_fsm/net210
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm__2286_ heichips25_can_lehmann_fsm/_1049_ heichips25_can_lehmann_fsm/net1209
+ heichips25_can_lehmann_fsm/_0599_ VPWR VGND sg13g2_xor2_1
XFILLER_0_505 VPWR VGND sg13g2_decap_8
XFILLER_0_527 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm_fanout298 heichips25_can_lehmann_fsm/net299 heichips25_can_lehmann_fsm/net298
+ VPWR VGND sg13g2_buf_1
Xclkbuf_2_2__f_clk clknet_2_2__leaf_clk clknet_0_clk VPWR VGND sg13g2_buf_16
XFILLER_28_277 VPWR VGND sg13g2_fill_1
XFILLER_11_122 VPWR VGND sg13g2_decap_4
XFILLER_24_483 VPWR VGND sg13g2_decap_8
XFILLER_24_494 VPWR VGND sg13g2_fill_1
XFILLER_40_976 VPWR VGND sg13g2_fill_1
XFILLER_11_177 VPWR VGND sg13g2_fill_1
XFILLER_22_62 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__1953_ VPWR heichips25_sap3/_1379_ heichips25_sap3__3965_/Q VGND
+ sg13g2_inv_1
XFILLER_22_95 VPWR VGND sg13g2_decap_8
XFILLER_4_877 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3623_ heichips25_sap3/_0124_ heichips25_sap3/_1111_ heichips25_sap3/_1183_
+ heichips25_sap3/net102 heichips25_sap3/_1403_ VPWR VGND sg13g2_a22oi_1
XFILLER_0_0 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3554_ heichips25_sap3__3959_/Q heichips25_sap3/_1138_ heichips25_sap3/_1134_
+ heichips25_sap3/_0100_ VPWR VGND sg13g2_mux2_1
Xheichips25_sap3__3485_ heichips25_sap3/_1083_ heichips25_sap3/_1081_ heichips25_sap3/_1082_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__2505_ heichips25_sap3/_1918_ heichips25_sap3/net88 heichips25_sap3__3948_/Q
+ heichips25_sap3/net89 heichips25_sap3__3940_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2436_ heichips25_sap3/_1734_ heichips25_sap3/_1846_ heichips25_sap3/_1849_
+ heichips25_sap3/_1850_ heichips25_sap3/_1851_ VPWR VGND sg13g2_and4_1
Xheichips25_sap3__2367_ heichips25_sap3/net256 heichips25_sap3/_1492_ heichips25_sap3/_1569_
+ heichips25_sap3/_1788_ VPWR VGND sg13g2_nor3_1
XFILLER_34_214 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2298_ heichips25_sap3/_1476_ heichips25_sap3/_1614_ heichips25_sap3/_1623_
+ heichips25_sap3/_1717_ heichips25_sap3/_1719_ VPWR VGND sg13g2_or4_1
XFILLER_16_973 VPWR VGND sg13g2_fill_1
XFILLER_31_921 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__4037_ heichips25_sap3/net460 VGND VPWR heichips25_sap3/net1012 heichips25_sap3__4037_/Q
+ clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_15_494 VPWR VGND sg13g2_decap_8
XFILLER_31_965 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2140_ heichips25_can_lehmann_fsm/_0479_ heichips25_can_lehmann_fsm/_0998_
+ heichips25_can_lehmann_fsm/_0477_ heichips25_can_lehmann_fsm/net315 heichips25_can_lehmann_fsm__2932_/Q
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2071_ VGND VPWR heichips25_can_lehmann_fsm/_0414_ heichips25_can_lehmann_fsm/_0415_
+ heichips25_can_lehmann_fsm/_0020_ heichips25_can_lehmann_fsm/_0416_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2973_ net732 VGND VPWR heichips25_can_lehmann_fsm/_0198_
+ heichips25_can_lehmann_fsm__2973_/Q clknet_leaf_6_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1924_ heichips25_can_lehmann_fsm/_1237_ heichips25_can_lehmann_fsm/net314
+ heichips25_can_lehmann_fsm__2936_/Q heichips25_can_lehmann_fsm/net318 heichips25_can_lehmann_fsm__3008_/Q
+ VPWR VGND sg13g2_a22oi_1
XFILLER_26_704 VPWR VGND sg13g2_fill_1
Xheichips25_sap3_fanout103 heichips25_sap3/_0767_ heichips25_sap3/net103 VPWR VGND
+ sg13g2_buf_1
Xheichips25_can_lehmann_fsm__1855_ heichips25_can_lehmann_fsm/_1168_ heichips25_can_lehmann_fsm/_1169_
+ heichips25_can_lehmann_fsm/_1167_ heichips25_can_lehmann_fsm/_1171_ VPWR VGND heichips25_can_lehmann_fsm/_1170_
+ sg13g2_nand4_1
Xheichips25_can_lehmann_fsm__2986__681 VPWR VGND net680 sg13g2_tiehi
Xheichips25_sap3_fanout114 heichips25_sap3/_0753_ heichips25_sap3/net114 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout125 heichips25_sap3/net126 heichips25_sap3/net125 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout136 heichips25_sap3/net137 heichips25_sap3/net136 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout147 heichips25_sap3/net149 heichips25_sap3/net147 VPWR VGND
+ sg13g2_buf_1
Xheichips25_can_lehmann_fsm__1786_ heichips25_can_lehmann_fsm/_0974_ heichips25_can_lehmann_fsm/_1100_
+ heichips25_can_lehmann_fsm/_1102_ VPWR VGND heichips25_can_lehmann_fsm/net1278 sg13g2_nand3b_1
Xheichips25_can_lehmann_fsm_hold1204 heichips25_can_lehmann_fsm/_0030_ VPWR VGND heichips25_can_lehmann_fsm/net1203
+ sg13g2_dlygate4sd3_1
Xheichips25_sap3_fanout169 heichips25_sap3/_1891_ heichips25_sap3/net169 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout158 heichips25_sap3/_0434_ heichips25_sap3/net158 VPWR VGND
+ sg13g2_buf_1
Xheichips25_can_lehmann_fsm_hold1215 heichips25_can_lehmann_fsm/_0288_ VPWR VGND heichips25_can_lehmann_fsm/net1214
+ sg13g2_dlygate4sd3_1
XFILLER_43_39 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm_hold1237 heichips25_can_lehmann_fsm__2806_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1236 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1248 heichips25_can_lehmann_fsm/_0014_ VPWR VGND heichips25_can_lehmann_fsm/net1247
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1259 heichips25_can_lehmann_fsm/_0007_ VPWR VGND heichips25_can_lehmann_fsm/net1258
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__2407_ VGND VPWR heichips25_can_lehmann_fsm/_0949_ heichips25_can_lehmann_fsm/net401
+ heichips25_can_lehmann_fsm/_0103_ heichips25_can_lehmann_fsm/_0669_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2338_ heichips25_can_lehmann_fsm/net474 VPWR heichips25_can_lehmann_fsm/_0635_
+ VGND heichips25_can_lehmann_fsm__2844_/Q heichips25_can_lehmann_fsm/net406 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2269_ heichips25_can_lehmann_fsm/net327 VPWR heichips25_can_lehmann_fsm/_0586_
+ VGND heichips25_can_lehmann_fsm/net1194 heichips25_can_lehmann_fsm/net207 sg13g2_o21ai_1
XFILLER_0_346 VPWR VGND sg13g2_decap_8
XFILLER_49_829 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3270_ heichips25_sap3/net123 heichips25_sap3/_0882_ heichips25_sap3/_0883_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__2221_ VGND VPWR heichips25_sap3/_1642_ heichips25_sap3/_1640_ heichips25_sap3/_1472_
+ sg13g2_or2_1
Xheichips25_can_lehmann_fsm__2965__765 VPWR VGND net764 sg13g2_tiehi
XFILLER_16_225 VPWR VGND sg13g2_decap_8
XFILLER_17_51 VPWR VGND sg13g2_decap_8
XFILLER_17_73 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2152_ heichips25_sap3/_1460_ heichips25_sap3/_1506_ heichips25_sap3/_1511_
+ heichips25_sap3/_1547_ heichips25_sap3/_1573_ VPWR VGND sg13g2_or4_1
XFILLER_31_206 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2083_ heichips25_sap3/_1437_ heichips25_sap3/_1438_ heichips25_sap3/net255
+ heichips25_sap3/_1501_ heichips25_sap3/_1504_ VPWR VGND sg13g2_or4_1
Xheichips25_can_lehmann_fsm__2861__774 VPWR VGND net773 sg13g2_tiehi
Xheichips25_sap3__2985_ heichips25_sap3/_0052_ heichips25_sap3/_0616_ heichips25_sap3/_0617_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__1936_ VPWR heichips25_sap3/_1362_ heichips25_sap3/net267 VGND sg13g2_inv_1
XFILLER_3_140 VPWR VGND sg13g2_decap_8
XFILLER_3_195 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3606_ heichips25_sap3/_1068_ heichips25_sap3__3974_/Q heichips25_sap3/net94
+ heichips25_sap3/_0115_ VPWR VGND sg13g2_mux2_1
Xheichips25_sap3__3537_ heichips25_sap3/_1127_ heichips25_sap3/_0888_ heichips25_sap3/_0870_
+ VPWR VGND sg13g2_nand2b_1
Xheichips25_sap3__3468_ heichips25_sap3/_0978_ heichips25_sap3/net121 net46 heichips25_sap3/_1069_
+ VPWR VGND sg13g2_a21o_1
Xheichips25_sap3__3399_ heichips25_sap3/net55 heichips25_sap3/_1005_ heichips25_sap3/_1006_
+ heichips25_sap3/_1007_ VPWR VGND sg13g2_nor3_1
Xheichips25_sap3__2419_ heichips25_sap3/_1836_ heichips25_sap3/_1834_ heichips25_sap3/_1835_
+ VPWR VGND sg13g2_nand2_1
XFILLER_35_545 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1640_ VPWR heichips25_can_lehmann_fsm/_0964_ heichips25_can_lehmann_fsm/net1002
+ VGND sg13g2_inv_1
XFILLER_22_217 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1571_ VPWR heichips25_can_lehmann_fsm/_0895_ heichips25_can_lehmann_fsm/net872
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__2907__682 VPWR VGND net681 sg13g2_tiehi
XFILLER_31_740 VPWR VGND sg13g2_decap_8
XFILLER_30_294 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2123_ VGND VPWR heichips25_can_lehmann_fsm__3024_/Q heichips25_can_lehmann_fsm/net312
+ heichips25_can_lehmann_fsm/_0462_ heichips25_can_lehmann_fsm/net303 sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2054_ heichips25_can_lehmann_fsm/_0402_ heichips25_can_lehmann_fsm/net347
+ heichips25_can_lehmann_fsm/net1255 VPWR VGND sg13g2_xnor2_1
X_20__522 VPWR VGND net521 sg13g2_tielo
Xheichips25_can_lehmann_fsm__2956_ net800 VGND VPWR heichips25_can_lehmann_fsm/_0181_
+ heichips25_can_lehmann_fsm__2956_/Q clknet_leaf_11_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1907_ heichips25_can_lehmann_fsm/_1220_ heichips25_can_lehmann_fsm/_0892_
+ heichips25_can_lehmann_fsm/net349 VPWR VGND sg13g2_nand2_1
Xheichips25_can_lehmann_fsm__2887_ net721 VGND VPWR heichips25_can_lehmann_fsm/_0112_
+ heichips25_can_lehmann_fsm__2887_/Q clknet_leaf_14_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1838_ heichips25_can_lehmann_fsm/_1154_ heichips25_can_lehmann_fsm__3059_/Q
+ heichips25_can_lehmann_fsm/net352 VPWR VGND sg13g2_xnor2_1
Xheichips25_can_lehmann_fsm_hold1001 heichips25_can_lehmann_fsm__2879_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1000 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__1769_ heichips25_can_lehmann_fsm/_1085_ heichips25_can_lehmann_fsm/net331
+ heichips25_can_lehmann_fsm__3038_/Q heichips25_can_lehmann_fsm/net317 heichips25_can_lehmann_fsm__2990_/Q
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm_hold1023 heichips25_can_lehmann_fsm__2981_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1022 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1056 heichips25_can_lehmann_fsm__2878_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1055 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1034 heichips25_can_lehmann_fsm__3018_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1033 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1045 heichips25_can_lehmann_fsm/_0280_ VPWR VGND heichips25_can_lehmann_fsm/net1044
+ sg13g2_dlygate4sd3_1
XFILLER_22_762 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm_hold1089 heichips25_can_lehmann_fsm__2841_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1088 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__2808__591 VPWR VGND net590 sg13g2_tiehi
Xheichips25_can_lehmann_fsm_hold1078 heichips25_can_lehmann_fsm__2951_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1077 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1067 heichips25_can_lehmann_fsm__2872_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1066 sg13g2_dlygate4sd3_1
XFILLER_21_272 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2839__529 VPWR VGND net528 sg13g2_tiehi
Xheichips25_sap3__2770_ heichips25_sap3/net169 heichips25_sap3/_1896_ heichips25_sap3/_0416_
+ VPWR VGND sg13g2_and2_1
XFILLER_0_121 VPWR VGND sg13g2_decap_8
XFILLER_1_699 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3322_ heichips25_sap3/_0865_ heichips25_sap3/_0888_ heichips25_sap3/_0853_
+ heichips25_sap3/_0933_ VPWR VGND sg13g2_nand3_1
XFILLER_29_372 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3253_ heichips25_sap3/_0866_ heichips25_sap3/net63 heichips25_sap3/_0820_
+ heichips25_sap3/_0864_ VPWR VGND sg13g2_and3_1
XFILLER_28_94 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3184_ heichips25_sap3/_0797_ heichips25_sap3/net132 heichips25_sap3__4000_/Q
+ heichips25_sap3/net139 heichips25_sap3__3984_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2204_ heichips25_sap3/_1625_ heichips25_sap3/_1546_ heichips25_sap3/_1566_
+ heichips25_sap3/_1477_ heichips25_sap3/_1463_ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2135_ heichips25_sap3/_1531_ VPWR heichips25_sap3/_1556_ VGND heichips25_sap3/_1545_
+ heichips25_sap3/_1555_ sg13g2_o21ai_1
XFILLER_40_581 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2066_ heichips25_sap3/net259 heichips25_sap3__3929_/Q heichips25_sap3/_1487_
+ VPWR VGND sg13g2_and2_1
XFILLER_5_43 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2968_ heichips25_sap3/_1767_ VPWR heichips25_sap3/_0605_ VGND heichips25_sap3/_0426_
+ heichips25_sap3/_0604_ sg13g2_o21ai_1
Xheichips25_sap3__2899_ heichips25_sap3/_0539_ heichips25_sap3/net159 heichips25_sap3/_0353_
+ VPWR VGND sg13g2_nand2b_1
Xheichips25_can_lehmann_fsm__2810_ net586 VGND VPWR heichips25_can_lehmann_fsm/_0035_
+ heichips25_can_lehmann_fsm__2810_/Q clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_27_309 VPWR VGND sg13g2_decap_8
XFILLER_47_180 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2741_ VGND VPWR heichips25_can_lehmann_fsm/_0860_ heichips25_can_lehmann_fsm/net391
+ heichips25_can_lehmann_fsm/_0270_ heichips25_can_lehmann_fsm/_0836_ sg13g2_a21oi_1
XFILLER_39_1015 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2672_ heichips25_can_lehmann_fsm/net482 VPWR heichips25_can_lehmann_fsm/_0802_
+ VGND heichips25_can_lehmann_fsm__3010_/Q heichips25_can_lehmann_fsm/net374 sg13g2_o21ai_1
XFILLER_23_504 VPWR VGND sg13g2_decap_8
XFILLER_35_386 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1623_ VPWR heichips25_can_lehmann_fsm/_0947_ heichips25_can_lehmann_fsm/net1000
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm_hold909 heichips25_can_lehmann_fsm__3041_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net908 sg13g2_dlygate4sd3_1
XFILLER_23_559 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2979__709 VPWR VGND net708 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__1554_ VPWR heichips25_can_lehmann_fsm/_0878_ heichips25_can_lehmann_fsm/net867
+ VGND sg13g2_inv_1
XFILLER_40_29 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2106_ VGND VPWR net18 heichips25_can_lehmann_fsm/net196
+ heichips25_can_lehmann_fsm/_0446_ heichips25_can_lehmann_fsm/net183 sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2037_ VPWR VGND heichips25_can_lehmann_fsm/net1227 heichips25_can_lehmann_fsm/net193
+ heichips25_can_lehmann_fsm/net189 heichips25_can_lehmann_fsm__2790_/Q heichips25_can_lehmann_fsm/_0387_
+ heichips25_can_lehmann_fsm/net198 sg13g2_a221oi_1
Xheichips25_can_lehmann_fsm__2939_ net579 VGND VPWR heichips25_can_lehmann_fsm/net1098
+ heichips25_can_lehmann_fsm__2939_/Q clknet_leaf_18_clk sg13g2_dfrbpq_1
XFILLER_26_331 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__3049__574 VPWR VGND net573 sg13g2_tiehi
XFILLER_26_353 VPWR VGND sg13g2_decap_4
XFILLER_27_876 VPWR VGND sg13g2_fill_1
XFILLER_42_857 VPWR VGND sg13g2_fill_1
XFILLER_42_824 VPWR VGND sg13g2_fill_1
XFILLER_41_323 VPWR VGND sg13g2_fill_2
XFILLER_26_386 VPWR VGND sg13g2_fill_1
XFILLER_26_397 VPWR VGND sg13g2_fill_1
XFILLER_10_743 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3940_ heichips25_sap3/net443 VGND VPWR heichips25_sap3/_0081_ heichips25_sap3__3940_/Q
+ heichips25_sap3__3988_/CLK sg13g2_dfrbpq_1
XFILLER_6_725 VPWR VGND sg13g2_fill_2
XFILLER_6_758 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2822_ heichips25_sap3/_0466_ heichips25_sap3/_0449_ heichips25_sap3/_0362_
+ heichips25_sap3/_0445_ heichips25_sap3/_0363_ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2753_ heichips25_sap3/_0399_ heichips25_sap3/_0350_ heichips25_sap3/_0397_
+ VPWR VGND sg13g2_xnor2_1
XFILLER_2_920 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2684_ heichips25_sap3/_0332_ VPWR heichips25_sap3/_0028_ VGND heichips25_sap3/_1382_
+ heichips25_sap3/net213 sg13g2_o21ai_1
XFILLER_2_986 VPWR VGND sg13g2_decap_8
XFILLER_37_629 VPWR VGND sg13g2_fill_1
XFILLER_37_618 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3305_ heichips25_sap3/_0916_ heichips25_sap3__3957_/Q heichips25_sap3/net145
+ VPWR VGND sg13g2_nand2_1
XFILLER_17_342 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3236_ heichips25_sap3/_0849_ heichips25_sap3/net133 heichips25_sap3__3996_/Q
+ heichips25_sap3/net140 heichips25_sap3__3988_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_17_397 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3167_ heichips25_sap3/_0780_ heichips25_sap3/net135 heichips25_sap3__3978_/Q
+ heichips25_sap3/net139 heichips25_sap3__3986_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_44_194 VPWR VGND sg13g2_decap_4
XFILLER_33_857 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2118_ heichips25_sap3/_1500_ heichips25_sap3/_1525_ heichips25_sap3/_1535_
+ heichips25_sap3/_1539_ VPWR VGND sg13g2_nor3_1
Xheichips25_sap3__3098_ heichips25_sap3/_1871_ VPWR heichips25_sap3/_0711_ VGND heichips25_sap3/net256
+ heichips25_sap3/_1569_ sg13g2_o21ai_1
Xheichips25_sap3__2049_ heichips25_sap3/_1454_ heichips25_sap3/net237 heichips25_sap3/_1470_
+ VPWR VGND sg13g2_nor2_1
XFILLER_4_290 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2724_ heichips25_can_lehmann_fsm/net479 VPWR heichips25_can_lehmann_fsm/_0828_
+ VGND heichips25_can_lehmann_fsm/net848 heichips25_can_lehmann_fsm/net410 sg13g2_o21ai_1
XFILLER_23_323 VPWR VGND sg13g2_decap_8
XFILLER_35_194 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2655_ VGND VPWR heichips25_can_lehmann_fsm/_0882_ heichips25_can_lehmann_fsm/net427
+ heichips25_can_lehmann_fsm/_0227_ heichips25_can_lehmann_fsm/_0793_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2586_ heichips25_can_lehmann_fsm/net476 VPWR heichips25_can_lehmann_fsm/_0759_
+ VGND heichips25_can_lehmann_fsm/net921 heichips25_can_lehmann_fsm/net396 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__1606_ VPWR heichips25_can_lehmann_fsm/_0930_ heichips25_can_lehmann_fsm/net909
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__1537_ VPWR heichips25_can_lehmann_fsm/_0861_ heichips25_can_lehmann_fsm/net877
+ VGND sg13g2_inv_1
XFILLER_15_824 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__4070_ heichips25_sap3__4070_/A uo_out_sap3\[1\] VPWR VGND sg13g2_buf_1
XFILLER_27_684 VPWR VGND sg13g2_decap_4
XFILLER_42_654 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3021_ VGND VPWR heichips25_sap3/_1365_ heichips25_sap3/net233 heichips25_sap3/_0069_
+ heichips25_sap3/_0636_ sg13g2_a21oi_1
XFILLER_26_183 VPWR VGND sg13g2_fill_2
XFILLER_14_389 VPWR VGND sg13g2_decap_8
XFILLER_6_500 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3923_ heichips25_sap3/net435 VGND VPWR heichips25_sap3/_0064_ heichips25_sap3__3923_/Q
+ clkload23/A sg13g2_dfrbpq_1
XFILLER_41_94 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3854_ VPWR VGND heichips25_sap3/_1348_ heichips25_sap3/_1353_ heichips25_sap3/_0286_
+ heichips25_sap3/_1359_ heichips25_sap3/_1354_ heichips25_sap3__4049_/Q sg13g2_a221oi_1
Xheichips25_sap3__2805_ heichips25_sap3/net159 VPWR heichips25_sap3/_0450_ VGND heichips25_sap3/net288
+ heichips25_sap3__3915_/Q sg13g2_o21ai_1
Xheichips25_sap3__3785_ heichips25_sap3/_1295_ heichips25_sap3/_1281_ heichips25_sap3__4013_/Q
+ heichips25_sap3/_1272_ heichips25_sap3__3973_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2736_ heichips25_sap3/_0380_ heichips25_sap3/_0381_ heichips25_sap3/_0350_
+ heichips25_sap3/_0382_ VPWR VGND sg13g2_nand3_1
XFILLER_2_772 VPWR VGND sg13g2_decap_8
XFILLER_49_231 VPWR VGND sg13g2_decap_8
XFILLER_38_905 VPWR VGND sg13g2_decap_8
XFILLER_2_11 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2667_ heichips25_sap3/net67 heichips25_sap3/_0247_ heichips25_sap3/_0256_
+ uio_oe_sap3\[2\] VPWR VGND sg13g2_nor3_1
XFILLER_49_275 VPWR VGND sg13g2_decap_8
XFILLER_38_927 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2598_ heichips25_sap3/net277 heichips25_sap3/net275 heichips25_sap3/_0270_
+ VPWR VGND sg13g2_xor2_1
XFILLER_18_695 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3219_ heichips25_sap3/_0717_ heichips25_sap3/net150 heichips25_sap3__4021_/Q
+ heichips25_sap3/_0832_ VPWR VGND sg13g2_nand3_1
XFILLER_33_643 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2440_ heichips25_can_lehmann_fsm/net464 VPWR heichips25_can_lehmann_fsm/_0686_
+ VGND heichips25_can_lehmann_fsm__2894_/Q heichips25_can_lehmann_fsm/net357 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2371_ VGND VPWR heichips25_can_lehmann_fsm/_0959_ heichips25_can_lehmann_fsm/net431
+ heichips25_can_lehmann_fsm/_0085_ heichips25_can_lehmann_fsm/_0651_ sg13g2_a21oi_1
XFILLER_20_348 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_fanout403 heichips25_can_lehmann_fsm/net408 heichips25_can_lehmann_fsm/net403
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout414 heichips25_can_lehmann_fsm/net420 heichips25_can_lehmann_fsm/net414
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout425 heichips25_can_lehmann_fsm/net432 heichips25_can_lehmann_fsm/net425
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout469 heichips25_can_lehmann_fsm/net470 heichips25_can_lehmann_fsm/net469
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm__3013__779 VPWR VGND net778 sg13g2_tiehi
XFILLER_28_448 VPWR VGND sg13g2_fill_1
XFILLER_37_960 VPWR VGND sg13g2_fill_1
XFILLER_37_982 VPWR VGND sg13g2_fill_1
XFILLER_23_131 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2707_ VGND VPWR heichips25_can_lehmann_fsm/_0868_ heichips25_can_lehmann_fsm/net384
+ heichips25_can_lehmann_fsm/_0253_ heichips25_can_lehmann_fsm/_0819_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2638_ heichips25_can_lehmann_fsm/net468 VPWR heichips25_can_lehmann_fsm/_0785_
+ VGND heichips25_can_lehmann_fsm/net1010 heichips25_can_lehmann_fsm/net398 sg13g2_o21ai_1
XFILLER_23_197 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2569_ VGND VPWR heichips25_can_lehmann_fsm/_0905_ heichips25_can_lehmann_fsm/net376
+ heichips25_can_lehmann_fsm/_0184_ heichips25_can_lehmann_fsm/_0750_ sg13g2_a21oi_1
XFILLER_3_525 VPWR VGND sg13g2_fill_2
XFILLER_2_4 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3570_ heichips25_sap3/_1097_ heichips25_sap3/_1149_ heichips25_sap3/_1150_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__2521_ heichips25_sap3/_1734_ heichips25_sap3/_1926_ heichips25_sap3/_1927_
+ heichips25_sap3/_1931_ heichips25_sap3/_0198_ VPWR VGND sg13g2_and4_1
XFILLER_47_713 VPWR VGND sg13g2_fill_1
XFILLER_47_702 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2452_ heichips25_sap3/_1447_ heichips25_sap3/net230 heichips25_sap3/net259
+ heichips25_sap3/_1865_ VPWR VGND sg13g2_nand3_1
XFILLER_47_735 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2383_ heichips25_sap3__3897_/Q net47 heichips25_sap3/net215 heichips25_sap3/_0038_
+ VPWR VGND sg13g2_mux2_1
XFILLER_28_960 VPWR VGND sg13g2_decap_8
XFILLER_46_278 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__4053_ heichips25_sap3/net453 VGND VPWR heichips25_sap3/net1144 heichips25_sap3__4053_/Q
+ clknet_leaf_22_clk sg13g2_dfrbpq_1
Xheichips25_sap3__3004_ heichips25_sap3__3919_/Q net46 heichips25_sap3/net202 heichips25_sap3/_0060_
+ VPWR VGND sg13g2_mux2_1
XFILLER_14_186 VPWR VGND sg13g2_decap_8
XFILLER_30_668 VPWR VGND sg13g2_fill_1
Xinput14 uio_in[3] net14 VPWR VGND sg13g2_buf_1
Xheichips25_sap3__3906_ heichips25_sap3/net455 VGND VPWR heichips25_sap3/_0047_ heichips25_sap3__3906_/Q
+ heichips25_sap3__3920_/CLK sg13g2_dfrbpq_1
XFILLER_6_385 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3837_ VPWR VGND heichips25_sap3/_1341_ heichips25_sap3/_0008_ heichips25_sap3/_1335_
+ heichips25_sap3/_1420_ heichips25_sap3/_1342_ heichips25_sap3/net291 sg13g2_a221oi_1
XFILLER_35_4 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3768_ heichips25_sap3/_1280_ heichips25_sap3/_1279_ heichips25_sap3__3963_/Q
+ heichips25_sap3/_1278_ heichips25_sap3__4003_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2719_ heichips25_sap3/_0364_ heichips25_sap3/_0363_ heichips25_sap3/_0362_
+ heichips25_sap3/_0365_ VPWR VGND sg13g2_a21o_1
Xheichips25_can_lehmann_fsm__2871__754 VPWR VGND net753 sg13g2_tiehi
Xheichips25_sap3__3699_ heichips25_sap3/_1232_ heichips25_sap3/net116 heichips25_sap3/_0876_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_can_lehmann_fsm__1940_ VGND VPWR heichips25_can_lehmann_fsm/_0293_ heichips25_can_lehmann_fsm/_0294_
+ heichips25_can_lehmann_fsm/_0303_ heichips25_can_lehmann_fsm/_0302_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__1871_ heichips25_can_lehmann_fsm/_1166_ heichips25_can_lehmann_fsm/net1172
+ heichips25_can_lehmann_fsm/_1185_ heichips25_can_lehmann_fsm/_1186_ VPWR VGND sg13g2_a21o_1
XFILLER_37_278 VPWR VGND sg13g2_decap_4
XFILLER_19_982 VPWR VGND sg13g2_fill_2
XFILLER_21_635 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2423_ VGND VPWR heichips25_can_lehmann_fsm/_0943_ heichips25_can_lehmann_fsm/net427
+ heichips25_can_lehmann_fsm/_0111_ heichips25_can_lehmann_fsm/_0677_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2354_ heichips25_can_lehmann_fsm/net495 VPWR heichips25_can_lehmann_fsm/_0643_
+ VGND heichips25_can_lehmann_fsm__2852_/Q heichips25_can_lehmann_fsm/net423 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2285_ VGND VPWR heichips25_can_lehmann_fsm/net207 heichips25_can_lehmann_fsm/_0597_
+ heichips25_can_lehmann_fsm/_0052_ heichips25_can_lehmann_fsm/_0598_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm_fanout200 heichips25_can_lehmann_fsm/_0305_ heichips25_can_lehmann_fsm/net200
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm__2917__662 VPWR VGND net661 sg13g2_tiehi
Xheichips25_can_lehmann_fsm_fanout299 heichips25_can_lehmann_fsm/_1002_ heichips25_can_lehmann_fsm/net299
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm__3048__606 VPWR VGND net605 sg13g2_tiehi
XFILLER_17_919 VPWR VGND sg13g2_decap_4
XFILLER_43_215 VPWR VGND sg13g2_decap_4
XFILLER_25_930 VPWR VGND sg13g2_decap_4
XFILLER_25_952 VPWR VGND sg13g2_fill_2
XFILLER_11_101 VPWR VGND sg13g2_decap_8
XFILLER_12_646 VPWR VGND sg13g2_decap_8
XFILLER_7_116 VPWR VGND sg13g2_fill_2
XFILLER_7_149 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__1952_ VPWR heichips25_sap3/_1378_ heichips25_sap3__3981_/Q VGND
+ sg13g2_inv_1
Xheichips25_sap3__3622_ heichips25_sap3/net102 heichips25_sap3/_0984_ heichips25_sap3/_1069_
+ heichips25_sap3/_1183_ VPWR VGND sg13g2_nor3_1
XFILLER_3_366 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2818__571 VPWR VGND net570 sg13g2_tiehi
Xheichips25_sap3__3553_ VGND VPWR heichips25_sap3/_1138_ heichips25_sap3/_1137_ heichips25_sap3/_1069_
+ sg13g2_or2_1
XFILLER_26_1028 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2504_ VPWR VGND heichips25_sap3__4020_/Q heichips25_sap3/net79 heichips25_sap3/net78
+ heichips25_sap3__4012_/Q heichips25_sap3/_1917_ heichips25_sap3/net218 sg13g2_a221oi_1
Xheichips25_sap3__3484_ VGND VPWR heichips25_sap3/net121 heichips25_sap3/_1045_ heichips25_sap3/_1082_
+ net47 sg13g2_a21oi_1
Xheichips25_sap3__2435_ heichips25_sap3/_1850_ heichips25_sap3/net73 heichips25_sap3__3999_/Q
+ heichips25_sap3/net77 heichips25_sap3__4015_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_35_727 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2366_ VGND VPWR heichips25_sap3/_1454_ heichips25_sap3/_1786_ heichips25_sap3/_1787_
+ heichips25_sap3/_1772_ sg13g2_a21oi_1
XFILLER_34_248 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2297_ heichips25_sap3/_1476_ heichips25_sap3/_1614_ heichips25_sap3/_1623_
+ heichips25_sap3/_1717_ heichips25_sap3/_1718_ VPWR VGND sg13g2_nor4_1
Xheichips25_sap3__4036_ heichips25_sap3/net461 VGND VPWR heichips25_sap3/net892 heichips25_sap3__4036_/Q
+ clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_8_32 VPWR VGND sg13g2_decap_8
XFILLER_8_65 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2899__698 VPWR VGND net697 sg13g2_tiehi
XFILLER_6_160 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2070_ heichips25_can_lehmann_fsm/net322 VPWR heichips25_can_lehmann_fsm/_0416_
+ VGND heichips25_can_lehmann_fsm/net347 heichips25_can_lehmann_fsm/net179 sg13g2_o21ai_1
XFILLER_38_521 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2972_ net736 VGND VPWR heichips25_can_lehmann_fsm/_0197_
+ heichips25_can_lehmann_fsm__2972_/Q clknet_leaf_14_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1923_ heichips25_can_lehmann_fsm/_1236_ heichips25_can_lehmann_fsm__2960_/Q
+ heichips25_can_lehmann_fsm/net307 VPWR VGND sg13g2_nand2_1
Xheichips25_sap3_rebuffer827 uio_out_sap3\[6\] heichips25_sap3/net826 VPWR VGND sg13g2_buf_1
Xheichips25_sap3_fanout104 heichips25_sap3/net105 heichips25_sap3/net104 VPWR VGND
+ sg13g2_buf_1
Xheichips25_can_lehmann_fsm__1854_ VGND VPWR heichips25_can_lehmann_fsm__2914_/Q heichips25_can_lehmann_fsm/net314
+ heichips25_can_lehmann_fsm/_1170_ heichips25_can_lehmann_fsm/net302 sg13g2_a21oi_1
X_19_ net520 uio_out_sap3\[5\] net504 net32 VPWR VGND sg13g2_mux2_1
Xheichips25_sap3_fanout126 heichips25_sap3/net130 heichips25_sap3/net126 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout115 heichips25_sap3/_0753_ heichips25_sap3/net115 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout137 heichips25_sap3/_0770_ heichips25_sap3/net137 VPWR VGND
+ sg13g2_buf_1
Xheichips25_can_lehmann_fsm__1785_ heichips25_can_lehmann_fsm/_1101_ heichips25_can_lehmann_fsm/_0974_
+ heichips25_can_lehmann_fsm/_1100_ VPWR VGND sg13g2_nand2_1
XFILLER_43_18 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm_hold1205 heichips25_can_lehmann_fsm__2834_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1204 sg13g2_dlygate4sd3_1
Xheichips25_sap3_fanout159 heichips25_sap3/_1895_ heichips25_sap3/net159 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout148 heichips25_sap3/net149 heichips25_sap3/net148 VPWR VGND
+ sg13g2_buf_1
Xheichips25_can_lehmann_fsm_hold1238 heichips25_can_lehmann_fsm/_0031_ VPWR VGND heichips25_can_lehmann_fsm/net1237
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1216 heichips25_can_lehmann_fsm__2804_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1215 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1227 heichips25_can_lehmann_fsm__2802_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1226 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1249 heichips25_can_lehmann_fsm__2783_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1248 sg13g2_dlygate4sd3_1
XFILLER_22_933 VPWR VGND sg13g2_fill_2
XFILLER_21_487 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2406_ heichips25_can_lehmann_fsm/net473 VPWR heichips25_can_lehmann_fsm/_0669_
+ VGND heichips25_can_lehmann_fsm/net1055 heichips25_can_lehmann_fsm/net401 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2337_ VGND VPWR heichips25_can_lehmann_fsm/_0967_ heichips25_can_lehmann_fsm/net367
+ heichips25_can_lehmann_fsm/_0068_ heichips25_can_lehmann_fsm/_0634_ sg13g2_a21oi_1
XFILLER_49_1028 VPWR VGND sg13g2_fill_1
XFILLER_49_1017 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2268_ VGND VPWR heichips25_can_lehmann_fsm/net941 heichips25_can_lehmann_fsm/net171
+ heichips25_can_lehmann_fsm/_0585_ heichips25_can_lehmann_fsm/_0584_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2199_ VPWR VGND heichips25_can_lehmann_fsm/_0530_ heichips25_can_lehmann_fsm/_1176_
+ heichips25_can_lehmann_fsm/_0529_ heichips25_can_lehmann_fsm/_0974_ heichips25_can_lehmann_fsm/_0034_
+ heichips25_can_lehmann_fsm/_0497_ sg13g2_a221oi_1
XFILLER_0_325 VPWR VGND sg13g2_decap_8
XFILLER_49_808 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2220_ heichips25_sap3/_1472_ heichips25_sap3/_1640_ heichips25_sap3/_1641_
+ VPWR VGND sg13g2_nor2_1
XFILLER_16_204 VPWR VGND sg13g2_decap_8
XFILLER_17_716 VPWR VGND sg13g2_fill_1
XFILLER_17_63 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2151_ heichips25_sap3/_1572_ heichips25_sap3/_1459_ heichips25_sap3/_1546_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__2082_ heichips25_sap3/_1437_ heichips25_sap3/_1438_ heichips25_sap3/net255
+ heichips25_sap3/_1501_ heichips25_sap3/_1503_ VPWR VGND sg13g2_nor4_1
XFILLER_8_458 VPWR VGND sg13g2_decap_8
XFILLER_12_498 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2984_ heichips25_sap3/_0617_ heichips25_sap3/net153 heichips25_sap3/_0406_
+ heichips25_sap3/net167 heichips25_sap3/net281 VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__1935_ VPWR heichips25_sap3/_1361_ heichips25_sap3/net260 VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__2972__737 VPWR VGND net736 sg13g2_tiehi
XFILLER_4_675 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3605_ heichips25_sap3/_1066_ heichips25_sap3__3973_/Q heichips25_sap3/net94
+ heichips25_sap3/_0114_ VPWR VGND sg13g2_mux2_1
Xheichips25_sap3__3536_ heichips25_sap3/_0094_ heichips25_sap3/_1124_ heichips25_sap3/_1126_
+ heichips25_sap3/net107 heichips25_sap3/_1418_ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3467_ heichips25_sap3/_1068_ heichips25_sap3__3942_/Q heichips25_sap3/net58
+ heichips25_sap3/_0083_ VPWR VGND sg13g2_mux2_1
XFILLER_12_6 VPWR VGND sg13g2_fill_1
XFILLER_35_513 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2418_ heichips25_sap3/_1835_ net8 heichips25_sap3/_1770_ VPWR VGND
+ sg13g2_nand2_1
Xheichips25_sap3__3398_ uio_out_sap3\[5\] heichips25_sap3/net828 heichips25_sap3/net68
+ heichips25_sap3/_1006_ VPWR VGND sg13g2_mux2_1
XFILLER_35_524 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2349_ heichips25_sap3/_1770_ heichips25_sap3/net231 heichips25_sap3/_1769_
+ VPWR VGND sg13g2_nand2_1
XFILLER_22_207 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1570_ VPWR heichips25_can_lehmann_fsm/_0894_ heichips25_can_lehmann_fsm/net1022
+ VGND sg13g2_inv_1
Xheichips25_sap3__4019_ heichips25_sap3/net456 VGND VPWR heichips25_sap3/_0160_ heichips25_sap3__4019_/Q
+ heichips25_sap3__4021_/CLK sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2122_ VPWR VGND heichips25_can_lehmann_fsm/_1163_ heichips25_can_lehmann_fsm/_0460_
+ heichips25_can_lehmann_fsm/_0453_ heichips25_can_lehmann_fsm__3047_/Q heichips25_can_lehmann_fsm/_0461_
+ heichips25_can_lehmann_fsm/_1166_ sg13g2_a221oi_1
Xheichips25_can_lehmann_fsm__2053_ heichips25_can_lehmann_fsm/_0401_ heichips25_can_lehmann_fsm/_0399_
+ heichips25_can_lehmann_fsm/_0400_ VPWR VGND sg13g2_xnor2_1
XFILLER_38_340 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2955_ net804 VGND VPWR heichips25_can_lehmann_fsm/net1028
+ heichips25_can_lehmann_fsm__2955_/Q clknet_leaf_11_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1906_ heichips25_can_lehmann_fsm/_1219_ heichips25_can_lehmann_fsm/net332
+ heichips25_can_lehmann_fsm__3057_/Q heichips25_can_lehmann_fsm/net314 heichips25_can_lehmann_fsm__2937_/Q
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2886_ net723 VGND VPWR heichips25_can_lehmann_fsm/net917
+ heichips25_can_lehmann_fsm__2886_/Q clknet_leaf_12_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1837_ heichips25_can_lehmann_fsm/_1153_ heichips25_can_lehmann_fsm/net348
+ heichips25_can_lehmann_fsm/_0996_ VPWR VGND sg13g2_nand2_1
XFILLER_41_527 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm_hold1002 heichips25_can_lehmann_fsm/_0105_ VPWR VGND heichips25_can_lehmann_fsm/net1001
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__1768_ VGND VPWR heichips25_can_lehmann_fsm/_1084_ heichips25_can_lehmann_fsm/net335
+ heichips25_can_lehmann_fsm__2870_/Q sg13g2_or2_1
Xheichips25_can_lehmann_fsm_hold1035 heichips25_can_lehmann_fsm__2846_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1034 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1046 heichips25_can_lehmann_fsm__2959_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1045 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1057 heichips25_can_lehmann_fsm__2899_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1056 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1024 heichips25_can_lehmann_fsm/_0206_ VPWR VGND heichips25_can_lehmann_fsm/net1023
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1079 heichips25_can_lehmann_fsm/_0176_ VPWR VGND heichips25_can_lehmann_fsm/net1078
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__1699_ heichips25_can_lehmann_fsm/_1023_ heichips25_can_lehmann_fsm/net294
+ heichips25_can_lehmann_fsm__2967_/Q heichips25_can_lehmann_fsm/net317 heichips25_can_lehmann_fsm__2991_/Q
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm_hold1068 heichips25_can_lehmann_fsm/_0098_ VPWR VGND heichips25_can_lehmann_fsm/net1067
+ sg13g2_dlygate4sd3_1
XFILLER_0_199 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3321_ heichips25_sap3/_0932_ heichips25_sap3/_0747_ heichips25_sap3/_0929_
+ heichips25_sap3/_0931_ VPWR VGND sg13g2_and3_1
XFILLER_28_84 VPWR VGND sg13g2_fill_2
XFILLER_29_351 VPWR VGND sg13g2_decap_8
XFILLER_17_546 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3252_ VGND VPWR heichips25_sap3/_0865_ heichips25_sap3/_0852_ heichips25_sap3/_0841_
+ sg13g2_or2_1
Xheichips25_sap3__3183_ heichips25_sap3/_0796_ heichips25_sap3/net148 heichips25_sap3__4008_/Q
+ heichips25_sap3/net116 heichips25_sap3__4024_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2203_ heichips25_sap3/_1624_ heichips25_sap3/net240 heichips25_sap3/_1623_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__2134_ heichips25_sap3/_1553_ VPWR heichips25_sap3/_1555_ VGND heichips25_sap3/_1460_
+ heichips25_sap3/_1552_ sg13g2_o21ai_1
XFILLER_12_251 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2065_ heichips25_sap3/_1486_ heichips25_sap3/_1477_ heichips25_sap3/_1468_
+ VPWR VGND sg13g2_nand2b_1
XFILLER_5_11 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2967_ heichips25_sap3/_0604_ heichips25_sap3/_1641_ heichips25_sap3/_1646_
+ VPWR VGND sg13g2_nand2_1
XFILLER_5_66 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2898_ uio_out_sap3\[5\] heichips25_sap3/net157 heichips25_sap3/_0538_
+ VPWR VGND sg13g2_nor2b_1
Xheichips25_sap3__3519_ heichips25_sap3/_1112_ heichips25_sap3/_1087_ uio_oe_sap3\[4\]
+ VPWR VGND sg13g2_nand2b_1
XFILLER_36_833 VPWR VGND sg13g2_fill_1
XFILLER_35_321 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2740_ heichips25_can_lehmann_fsm/net470 VPWR heichips25_can_lehmann_fsm/_0836_
+ VGND heichips25_can_lehmann_fsm/net1154 heichips25_can_lehmann_fsm/net391 sg13g2_o21ai_1
XFILLER_39_1027 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2671_ VGND VPWR heichips25_can_lehmann_fsm/_0878_ heichips25_can_lehmann_fsm/net416
+ heichips25_can_lehmann_fsm/_0235_ heichips25_can_lehmann_fsm/_0801_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__1622_ VPWR heichips25_can_lehmann_fsm/_0946_ heichips25_can_lehmann_fsm/net1095
+ VGND sg13g2_inv_1
XFILLER_23_527 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__1553_ VPWR heichips25_can_lehmann_fsm/_0877_ heichips25_can_lehmann_fsm/net881
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__2105_ heichips25_can_lehmann_fsm/_0444_ heichips25_can_lehmann_fsm/_0441_
+ heichips25_can_lehmann_fsm/net196 heichips25_can_lehmann_fsm/_0445_ VPWR VGND sg13g2_a21o_1
Xheichips25_can_lehmann_fsm__3016__755 VPWR VGND net754 sg13g2_tiehi
XFILLER_49_39 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2036_ heichips25_can_lehmann_fsm__2783_/Q heichips25_can_lehmann_fsm/net193
+ heichips25_can_lehmann_fsm/_0386_ VPWR VGND sg13g2_nor2b_1
XFILLER_27_811 VPWR VGND sg13g2_fill_2
XFILLER_38_181 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2938_ net583 VGND VPWR heichips25_can_lehmann_fsm/net1014
+ heichips25_can_lehmann_fsm__2938_/Q clknet_leaf_17_clk sg13g2_dfrbpq_1
XFILLER_27_822 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2869_ net757 VGND VPWR heichips25_can_lehmann_fsm/net988
+ heichips25_can_lehmann_fsm__2869_/Q clknet_leaf_20_clk sg13g2_dfrbpq_1
XFILLER_26_365 VPWR VGND sg13g2_decap_8
XFILLER_14_549 VPWR VGND sg13g2_decap_8
XFILLER_14_31 VPWR VGND sg13g2_fill_2
XFILLER_5_203 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3870_ heichips25_sap3__3889_/Q heichips25_sap3/net1112 heichips25_sap3/net341
+ heichips25_sap3/_0197_ VPWR VGND sg13g2_mux2_1
XFILLER_10_777 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2821_ VPWR VGND heichips25_sap3/net289 heichips25_sap3/_0464_ heichips25_sap3/_0417_
+ heichips25_sap3/net285 heichips25_sap3/_0465_ heichips25_sap3/_0416_ sg13g2_a221oi_1
XFILLER_5_258 VPWR VGND sg13g2_fill_1
XFILLER_5_247 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2752_ heichips25_sap3/_0350_ heichips25_sap3/_0397_ heichips25_sap3/_0398_
+ VPWR VGND sg13g2_nor2b_1
Xheichips25_sap3__2683_ heichips25_sap3/_0332_ heichips25_sap3__3887_/Q heichips25_sap3/net213
+ VPWR VGND sg13g2_nand2_1
XFILLER_2_965 VPWR VGND sg13g2_decap_8
XFILLER_18_844 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3304_ VPWR VGND heichips25_sap3__3997_/Q heichips25_sap3/net128
+ heichips25_sap3/net147 heichips25_sap3__4013_/Q heichips25_sap3/_0915_ heichips25_sap3/net116
+ sg13g2_a221oi_1
XFILLER_45_663 VPWR VGND sg13g2_fill_2
XFILLER_17_354 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3235_ heichips25_sap3/_0848_ heichips25_sap3/net138 heichips25_sap3__3980_/Q
+ heichips25_sap3/net145 heichips25_sap3__3964_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__3028__659 VPWR VGND net658 sg13g2_tiehi
XFILLER_45_674 VPWR VGND sg13g2_fill_2
XFILLER_32_313 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3166_ heichips25_sap3/_0779_ heichips25_sap3/net147 heichips25_sap3__4010_/Q
+ heichips25_sap3/net117 heichips25_sap3__4026_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_32_357 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3097_ VGND VPWR heichips25_sap3/_1510_ heichips25_sap3/_0708_ heichips25_sap3/_0710_
+ heichips25_sap3/net222 sg13g2_a21oi_1
Xheichips25_sap3__2117_ heichips25_sap3/_1525_ heichips25_sap3/_1535_ heichips25_sap3/_1538_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__2048_ VPWR VGND heichips25_sap3/net247 heichips25_sap3/_1455_ heichips25_sap3/_1468_
+ heichips25_sap3/net249 heichips25_sap3/_1469_ heichips25_sap3/net234 sg13g2_a221oi_1
XFILLER_9_564 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3999_ heichips25_sap3/net438 VGND VPWR heichips25_sap3/_0140_ heichips25_sap3__3999_/Q
+ heichips25_sap3__4017_/CLK sg13g2_dfrbpq_1
XFILLER_5_781 VPWR VGND sg13g2_decap_8
XFILLER_45_1020 VPWR VGND sg13g2_decap_8
XFILLER_28_619 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2723_ VGND VPWR heichips25_can_lehmann_fsm/_0864_ heichips25_can_lehmann_fsm/net369
+ heichips25_can_lehmann_fsm/_0261_ heichips25_can_lehmann_fsm/_0827_ sg13g2_a21oi_1
XFILLER_24_803 VPWR VGND sg13g2_decap_4
XFILLER_24_814 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2881__734 VPWR VGND net733 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2654_ heichips25_can_lehmann_fsm/net497 VPWR heichips25_can_lehmann_fsm/_0793_
+ VGND heichips25_can_lehmann_fsm/net1134 heichips25_can_lehmann_fsm/net427 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2585_ VGND VPWR heichips25_can_lehmann_fsm/_0901_ heichips25_can_lehmann_fsm/net358
+ heichips25_can_lehmann_fsm/_0192_ heichips25_can_lehmann_fsm/_0758_ sg13g2_a21oi_1
XFILLER_11_519 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1605_ VPWR heichips25_can_lehmann_fsm/_0929_ heichips25_can_lehmann_fsm/net966
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__1536_ VPWR heichips25_can_lehmann_fsm/_0860_ heichips25_can_lehmann_fsm/net1229
+ VGND sg13g2_inv_1
XFILLER_3_729 VPWR VGND sg13g2_fill_2
XFILLER_2_239 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2019_ heichips25_can_lehmann_fsm/net321 VPWR heichips25_can_lehmann_fsm/_0372_
+ VGND heichips25_can_lehmann_fsm/net1259 heichips25_can_lehmann_fsm/net178 sg13g2_o21ai_1
Xheichips25_sap3__3020_ heichips25_sap3/net233 uio_out_sap3\[5\] heichips25_sap3/_0636_
+ VPWR VGND sg13g2_nor2_1
XFILLER_41_132 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2782__643 VPWR VGND net642 sg13g2_tiehi
XFILLER_30_839 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2997__618 VPWR VGND net617 sg13g2_tiehi
XFILLER_6_545 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3922_ heichips25_sap3/net450 VGND VPWR heichips25_sap3/_0063_ heichips25_sap3__3922_/Q
+ heichips25_sap3__3922_/CLK sg13g2_dfrbpq_1
Xheichips25_sap3__3853_ heichips25_sap3/_1353_ heichips25_sap3__4058_/Q heichips25_sap3__4048_/Q
+ heichips25_sap3/_1352_ VPWR VGND sg13g2_and3_1
Xheichips25_sap3__2804_ heichips25_sap3/_1885_ heichips25_sap3/net169 heichips25_sap3/_0449_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__3784_ heichips25_sap3/net339 heichips25_sap3/net1141 heichips25_sap3/_1294_
+ heichips25_sap3/_0174_ VPWR VGND sg13g2_a21o_1
Xheichips25_sap3__2735_ heichips25_sap3/_0347_ heichips25_sap3/_0348_ heichips25_sap3/_0381_
+ VPWR VGND sg13g2_nor2b_1
XFILLER_29_1026 VPWR VGND sg13g2_fill_2
XFILLER_2_784 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2666_ VPWR heichips25_sap3/_0327_ uio_oe_sap3\[1\] VGND sg13g2_inv_1
XFILLER_2_67 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2597_ heichips25_sap3/_0269_ heichips25_sap3/_1801_ net44 VPWR VGND
+ sg13g2_nand2_1
XFILLER_2_78 VPWR VGND sg13g2_fill_1
XFILLER_2_89 VPWR VGND sg13g2_fill_1
XFILLER_18_674 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2828__551 VPWR VGND net550 sg13g2_tiehi
XFILLER_17_184 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3218_ heichips25_sap3/_0831_ heichips25_sap3__4005_/Q heichips25_sap3/net147
+ VPWR VGND sg13g2_nand2_1
XFILLER_32_121 VPWR VGND sg13g2_decap_8
XFILLER_33_633 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3149_ heichips25_sap3/_0666_ heichips25_sap3/_0678_ heichips25_sap3/_0762_
+ VPWR VGND sg13g2_nor2_1
XFILLER_33_688 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2370_ heichips25_can_lehmann_fsm/net501 VPWR heichips25_can_lehmann_fsm/_0651_
+ VGND heichips25_can_lehmann_fsm/net980 heichips25_can_lehmann_fsm/net431 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm_fanout404 heichips25_can_lehmann_fsm/net405 heichips25_can_lehmann_fsm/net404
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout415 heichips25_can_lehmann_fsm/net416 heichips25_can_lehmann_fsm/net415
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout426 heichips25_can_lehmann_fsm/net429 heichips25_can_lehmann_fsm/net426
+ VPWR VGND sg13g2_buf_1
XFILLER_37_972 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2706_ heichips25_can_lehmann_fsm/net502 VPWR heichips25_can_lehmann_fsm/_0819_
+ VGND heichips25_can_lehmann_fsm/net1153 heichips25_can_lehmann_fsm/net385 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2637_ VGND VPWR heichips25_can_lehmann_fsm/_0888_ heichips25_can_lehmann_fsm/net357
+ heichips25_can_lehmann_fsm/_0218_ heichips25_can_lehmann_fsm/_0784_ sg13g2_a21oi_1
XFILLER_24_666 VPWR VGND sg13g2_decap_4
XFILLER_12_839 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2568_ heichips25_can_lehmann_fsm/net487 VPWR heichips25_can_lehmann_fsm/_0750_
+ VGND heichips25_can_lehmann_fsm/net1109 heichips25_can_lehmann_fsm/net376 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2499_ VGND VPWR heichips25_can_lehmann_fsm/_0923_ heichips25_can_lehmann_fsm/net391
+ heichips25_can_lehmann_fsm/_0149_ heichips25_can_lehmann_fsm/_0715_ sg13g2_a21oi_1
XFILLER_11_54 VPWR VGND sg13g2_decap_8
XFILLER_11_65 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2520_ heichips25_sap3/_1931_ heichips25_sap3/net74 heichips25_sap3__3995_/Q
+ heichips25_sap3/net78 heichips25_sap3__4011_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2451_ heichips25_sap3__3894_/Q net46 heichips25_sap3/net215 heichips25_sap3/_0035_
+ VPWR VGND sg13g2_mux2_1
Xheichips25_sap3__2382_ heichips25_sap3/_1494_ heichips25_sap3/net227 heichips25_sap3/_1441_
+ heichips25_sap3/_1802_ VPWR VGND sg13g2_nand3_1
Xheichips25_can_lehmann_fsm__2968__753 VPWR VGND net752 sg13g2_tiehi
Xheichips25_sap3__4052_ heichips25_sap3/net452 VGND VPWR heichips25_sap3/_0193_ heichips25_sap3__4052_/Q
+ clknet_leaf_23_clk sg13g2_dfrbpq_1
XFILLER_15_633 VPWR VGND sg13g2_decap_8
XFILLER_14_143 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3003_ VGND VPWR heichips25_sap3/net45 heichips25_sap3/net201 heichips25_sap3/_0059_
+ heichips25_sap3/_0628_ sg13g2_a21oi_1
XFILLER_14_165 VPWR VGND sg13g2_decap_8
Xinput15 uio_in[4] net15 VPWR VGND sg13g2_buf_1
XFILLER_7_854 VPWR VGND sg13g2_fill_1
XFILLER_6_331 VPWR VGND sg13g2_fill_2
XFILLER_10_393 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3905_ heichips25_sap3/net455 VGND VPWR heichips25_sap3/_0046_ heichips25_sap3__3905_/Q
+ clkload26/A sg13g2_dfrbpq_1
Xheichips25_sap3__3836_ VPWR VGND heichips25_sap3__3954_/Q heichips25_sap3/_1340_
+ heichips25_sap3/_1282_ heichips25_sap3__4018_/Q heichips25_sap3/_1341_ heichips25_sap3/_1281_
+ sg13g2_a221oi_1
Xheichips25_sap3__3767_ heichips25_sap3__4040_/Q heichips25_sap3__4041_/Q heichips25_sap3/_1257_
+ heichips25_sap3/_1279_ VPWR VGND sg13g2_nor3_1
Xheichips25_sap3__2718_ heichips25_sap3/net288 heichips25_sap3__3915_/Q heichips25_sap3/_0364_
+ VPWR VGND sg13g2_and2_1
Xheichips25_sap3__3698_ heichips25_sap3/_1231_ heichips25_sap3__4011_/Q heichips25_sap3/net115
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__2649_ heichips25_sap3/net224 heichips25_sap3/_0315_ heichips25_sap3/_1480_
+ heichips25_sap3/_0316_ VPWR VGND sg13g2_nand3_1
XFILLER_38_736 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1870_ heichips25_can_lehmann_fsm/_1184_ VPWR heichips25_can_lehmann_fsm/_1185_
+ VGND heichips25_can_lehmann_fsm/net219 heichips25_can_lehmann_fsm/_1183_ sg13g2_o21ai_1
XFILLER_46_791 VPWR VGND sg13g2_fill_2
XFILLER_34_931 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2422_ heichips25_can_lehmann_fsm/net498 VPWR heichips25_can_lehmann_fsm/_0677_
+ VGND heichips25_can_lehmann_fsm__2886_/Q heichips25_can_lehmann_fsm/net427 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2353_ VGND VPWR heichips25_can_lehmann_fsm/_0963_ heichips25_can_lehmann_fsm/net383
+ heichips25_can_lehmann_fsm/_0076_ heichips25_can_lehmann_fsm/_0642_ sg13g2_a21oi_1
Xclkbuf_leaf_9_clk clknet_2_3__leaf_clk clknet_leaf_9_clk VPWR VGND sg13g2_buf_8
Xheichips25_can_lehmann_fsm__2284_ heichips25_can_lehmann_fsm/net328 VPWR heichips25_can_lehmann_fsm/_0598_
+ VGND heichips25_can_lehmann_fsm/net1170 heichips25_can_lehmann_fsm/net207 sg13g2_o21ai_1
XFILLER_28_213 VPWR VGND sg13g2_decap_8
XFILLER_43_205 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__1999_ heichips25_can_lehmann_fsm/_0354_ heichips25_can_lehmann_fsm/_0352_
+ heichips25_can_lehmann_fsm/_0353_ heichips25_can_lehmann_fsm/_0355_ VPWR VGND sg13g2_a21o_1
XFILLER_16_419 VPWR VGND sg13g2_fill_1
XFILLER_40_989 VPWR VGND sg13g2_fill_1
XFILLER_12_658 VPWR VGND sg13g2_fill_1
XFILLER_11_168 VPWR VGND sg13g2_decap_4
XFILLER_22_42 VPWR VGND sg13g2_fill_2
XFILLER_22_53 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__1951_ VPWR heichips25_sap3/_1377_ heichips25_sap3__3997_/Q VGND
+ sg13g2_inv_1
XFILLER_3_334 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3621_ heichips25_sap3/_0123_ heichips25_sap3/_1106_ heichips25_sap3/_1182_
+ heichips25_sap3/net102 heichips25_sap3/_1371_ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3552_ heichips25_sap3/net99 heichips25_sap3/_0973_ heichips25_sap3/_1137_
+ VPWR VGND sg13g2_and2_1
Xheichips25_sap3__2503_ heichips25_sap3/_1914_ heichips25_sap3/_1915_ heichips25_sap3/_1916_
+ VPWR VGND sg13g2_and2_1
XFILLER_47_500 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3483_ heichips25_sap3/_1081_ heichips25_sap3/net98 heichips25_sap3/_1038_
+ VPWR VGND sg13g2_nand2_1
XFILLER_19_213 VPWR VGND sg13g2_decap_4
XFILLER_47_83 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2434_ heichips25_sap3/_1849_ heichips25_sap3/net72 heichips25_sap3__3975_/Q
+ heichips25_sap3/net217 heichips25_sap3__4007_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_19_235 VPWR VGND sg13g2_decap_8
XFILLER_19_246 VPWR VGND sg13g2_fill_1
XFILLER_47_588 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2365_ VGND VPWR heichips25_sap3/_1641_ heichips25_sap3/_1781_ heichips25_sap3/_1786_
+ heichips25_sap3/_1785_ sg13g2_a21oi_1
XFILLER_19_279 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2296_ heichips25_sap3/_1435_ heichips25_sap3/_1613_ heichips25_sap3/_1717_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__4035_ heichips25_sap3/net458 VGND VPWR heichips25_sap3/net926 heichips25_sap3__4035_/Q
+ clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_42_282 VPWR VGND sg13g2_decap_8
XFILLER_42_271 VPWR VGND sg13g2_fill_2
XFILLER_8_11 VPWR VGND sg13g2_decap_4
XFILLER_8_99 VPWR VGND sg13g2_decap_8
XFILLER_8_88 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm_hold890 heichips25_can_lehmann_fsm__2987_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net889 sg13g2_dlygate4sd3_1
XFILLER_6_194 VPWR VGND sg13g2_fill_2
XFILLER_6_183 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3819_ VPWR VGND heichips25_sap3/_1325_ heichips25_sap3/net340 heichips25_sap3/_1319_
+ heichips25_sap3/_1404_ heichips25_sap3/_1326_ heichips25_sap3/net291 sg13g2_a221oi_1
Xclkbuf_5_10__f_heichips25_sap3\_sap_3_inst.alu_inst.clk heichips25_sap3__4016_/CLK
+ clknet_4_5_0_heichips25_sap3\/sap_3_inst.alu_inst.clk VPWR VGND sg13g2_buf_16
XFILLER_38_511 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2971_ net740 VGND VPWR heichips25_can_lehmann_fsm/net947
+ heichips25_can_lehmann_fsm__2971_/Q clknet_leaf_21_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1922_ heichips25_can_lehmann_fsm/_1224_ heichips25_can_lehmann_fsm/_1223_
+ heichips25_can_lehmann_fsm/_1233_ heichips25_can_lehmann_fsm/_1235_ VPWR VGND sg13g2_a21o_1
XFILLER_38_577 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1853_ heichips25_can_lehmann_fsm/_1169_ heichips25_can_lehmann_fsm/net295
+ heichips25_can_lehmann_fsm__2962_/Q heichips25_can_lehmann_fsm/net332 heichips25_can_lehmann_fsm__3034_/Q
+ VPWR VGND sg13g2_a22oi_1
X_18_ net519 net46 net504 net31 VPWR VGND sg13g2_mux2_1
Xheichips25_sap3_fanout105 heichips25_sap3/_0763_ heichips25_sap3/net105 VPWR VGND
+ sg13g2_buf_1
XFILLER_26_728 VPWR VGND sg13g2_decap_4
Xheichips25_sap3_fanout116 heichips25_sap3/net118 heichips25_sap3/net116 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout138 heichips25_sap3/net139 heichips25_sap3/net138 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_rebuffer828 heichips25_sap3/_1736_ heichips25_sap3/net827 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout127 heichips25_sap3/net130 heichips25_sap3/net127 VPWR VGND
+ sg13g2_buf_1
XFILLER_25_227 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1784_ heichips25_can_lehmann_fsm/net1192 heichips25_can_lehmann_fsm__2807_/Q
+ heichips25_can_lehmann_fsm__2806_/Q heichips25_can_lehmann_fsm/_1098_ heichips25_can_lehmann_fsm/_1100_
+ VPWR VGND sg13g2_nor4_1
Xheichips25_can_lehmann_fsm_hold1206 heichips25_can_lehmann_fsm__2817_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1205 sg13g2_dlygate4sd3_1
Xheichips25_sap3_fanout149 heichips25_sap3/_0754_ heichips25_sap3/net149 VPWR VGND
+ sg13g2_buf_1
Xheichips25_can_lehmann_fsm_hold1217 heichips25_can_lehmann_fsm/_0029_ VPWR VGND heichips25_can_lehmann_fsm/net1216
+ sg13g2_dlygate4sd3_1
XFILLER_40_219 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_hold1228 heichips25_can_lehmann_fsm__2792_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1227 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1239 heichips25_can_lehmann_fsm__2791_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1238 sg13g2_dlygate4sd3_1
Xheichips25_sap3_hold926 heichips25_sap3__4035_/Q VPWR VGND heichips25_sap3/net925
+ sg13g2_dlygate4sd3_1
XFILLER_22_989 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2405_ VGND VPWR heichips25_can_lehmann_fsm/_0950_ heichips25_can_lehmann_fsm/net401
+ heichips25_can_lehmann_fsm/_0102_ heichips25_can_lehmann_fsm/_0668_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2336_ heichips25_can_lehmann_fsm/net474 VPWR heichips25_can_lehmann_fsm/_0634_
+ VGND heichips25_can_lehmann_fsm/net974 heichips25_can_lehmann_fsm/net364 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__3019__731 VPWR VGND net730 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2267_ heichips25_can_lehmann_fsm/net171 heichips25_can_lehmann_fsm/_0583_
+ heichips25_can_lehmann_fsm/_0584_ VPWR VGND sg13g2_nor2_1
Xheichips25_can_lehmann_fsm__2198_ VPWR VGND net18 heichips25_can_lehmann_fsm/_0497_
+ heichips25_can_lehmann_fsm/_0499_ heichips25_can_lehmann_fsm/net1088 heichips25_can_lehmann_fsm/_0530_
+ heichips25_can_lehmann_fsm/net175 sg13g2_a221oi_1
XFILLER_0_304 VPWR VGND sg13g2_decap_8
XFILLER_29_577 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2150_ VGND VPWR heichips25_sap3/_1544_ heichips25_sap3/_1570_ heichips25_sap3/_1571_
+ heichips25_sap3/_1565_ sg13g2_a21oi_1
XFILLER_44_569 VPWR VGND sg13g2_decap_8
XFILLER_17_75 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2081_ heichips25_sap3/_1437_ heichips25_sap3/_1501_ heichips25_sap3/_1502_
+ VPWR VGND sg13g2_nor2_1
XFILLER_25_783 VPWR VGND sg13g2_decap_4
XFILLER_12_444 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2983_ heichips25_sap3/_0616_ heichips25_sap3__3911_/Q heichips25_sap3/_0607_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__1934_ VPWR heichips25_sap3/_1360_ heichips25_sap3/net1130 VGND sg13g2_inv_1
XFILLER_3_175 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3604_ heichips25_sap3/_1175_ heichips25_sap3__3972_/Q heichips25_sap3/net94
+ heichips25_sap3/_0113_ VPWR VGND sg13g2_mux2_1
Xheichips25_sap3__3535_ heichips25_sap3/net107 heichips25_sap3/_1125_ heichips25_sap3/_1126_
+ VPWR VGND sg13g2_nor2_1
XFILLER_48_853 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3466_ heichips25_sap3/_0947_ heichips25_sap3/net98 heichips25_sap3/_1067_
+ heichips25_sap3/_1068_ VPWR VGND sg13g2_a21o_1
Xheichips25_sap3__2417_ heichips25_sap3/_1833_ VPWR heichips25_sap3/_1834_ VGND heichips25_sap3/net279
+ heichips25_sap3/net155 sg13g2_o21ai_1
Xheichips25_sap3__3397_ VGND VPWR heichips25_sap3/net124 heichips25_sap3/_1001_ heichips25_sap3/_1005_
+ heichips25_sap3/_1004_ sg13g2_a21oi_1
Xheichips25_sap3__2348_ heichips25_sap3/_1769_ heichips25_sap3/_1753_ heichips25_sap3/_1768_
+ VPWR VGND sg13g2_nand2_1
XFILLER_16_761 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2279_ heichips25_sap3/_1659_ heichips25_sap3/_1660_ heichips25_sap3/_1698_
+ heichips25_sap3/_1699_ heichips25_sap3/_1700_ VPWR VGND sg13g2_and4_1
XFILLER_15_260 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__4018_ heichips25_sap3/net442 VGND VPWR heichips25_sap3/_0159_ heichips25_sap3__4018_/Q
+ heichips25_sap3__4018_/CLK sg13g2_dfrbpq_1
XFILLER_30_230 VPWR VGND sg13g2_fill_1
XFILLER_30_274 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2121_ heichips25_can_lehmann_fsm/_1090_ VPWR heichips25_can_lehmann_fsm/_0460_
+ VGND heichips25_can_lehmann_fsm/net219 heichips25_can_lehmann_fsm/_0459_ sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2052_ heichips25_can_lehmann_fsm/net344 heichips25_can_lehmann_fsm__2801_/Q
+ heichips25_can_lehmann_fsm/_0400_ VPWR VGND sg13g2_xor2_1
Xheichips25_can_lehmann_fsm__2954_ net808 VGND VPWR heichips25_can_lehmann_fsm/net1104
+ heichips25_can_lehmann_fsm__2954_/Q clknet_leaf_10_clk sg13g2_dfrbpq_1
XFILLER_39_864 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1905_ heichips25_can_lehmann_fsm/_1218_ heichips25_can_lehmann_fsm/net307
+ heichips25_can_lehmann_fsm__2961_/Q heichips25_can_lehmann_fsm/net311 heichips25_can_lehmann_fsm__3033_/Q
+ VPWR VGND sg13g2_a22oi_1
XFILLER_26_503 VPWR VGND sg13g2_fill_1
XFILLER_0_1020 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2885_ net725 VGND VPWR heichips25_can_lehmann_fsm/_0110_
+ heichips25_can_lehmann_fsm__2885_/Q clknet_leaf_12_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1836_ heichips25_can_lehmann_fsm/_1151_ VPWR heichips25_can_lehmann_fsm/_1152_
+ VGND heichips25_can_lehmann_fsm/_1074_ heichips25_can_lehmann_fsm/_1144_ sg13g2_o21ai_1
XFILLER_41_539 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm_hold1003 heichips25_can_lehmann_fsm__2849_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1002 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1014 heichips25_can_lehmann_fsm__2937_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1013 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__1767_ uo_out_fsm\[7\] heichips25_can_lehmann_fsm/_1082_
+ heichips25_can_lehmann_fsm/_1083_ VPWR VGND sg13g2_nand2_1
Xheichips25_can_lehmann_fsm_hold1025 heichips25_can_lehmann_fsm__2902_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1024 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1047 heichips25_can_lehmann_fsm/_0185_ VPWR VGND heichips25_can_lehmann_fsm/net1046
+ sg13g2_dlygate4sd3_1
XFILLER_21_230 VPWR VGND sg13g2_decap_4
XFILLER_22_742 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_hold1036 heichips25_can_lehmann_fsm__2957_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1035 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1069 heichips25_can_lehmann_fsm__2868_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1068 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__1698_ heichips25_can_lehmann_fsm/_1021_ VPWR heichips25_can_lehmann_fsm/_1022_
+ VGND heichips25_can_lehmann_fsm__2872_/Q heichips25_can_lehmann_fsm/net336 sg13g2_o21ai_1
XFILLER_16_1028 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_hold1058 heichips25_can_lehmann_fsm/_0124_ VPWR VGND heichips25_can_lehmann_fsm/net1057
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__2319_ VGND VPWR heichips25_can_lehmann_fsm/_0972_ heichips25_can_lehmann_fsm/net401
+ heichips25_can_lehmann_fsm/_0059_ heichips25_can_lehmann_fsm/_0625_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2891__714 VPWR VGND net713 sg13g2_tiehi
XFILLER_0_112 VPWR VGND sg13g2_decap_4
XFILLER_0_178 VPWR VGND sg13g2_fill_2
XFILLER_0_167 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3320_ heichips25_sap3/_0930_ VPWR heichips25_sap3/_0931_ VGND net44
+ heichips25_sap3/net68 sg13g2_o21ai_1
Xheichips25_sap3__3251_ heichips25_sap3/_0864_ heichips25_sap3/_0850_ heichips25_sap3/_0851_
+ heichips25_sap3/_0840_ heichips25_sap3/_0835_ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2202_ heichips25_sap3/_1448_ heichips25_sap3/_1488_ heichips25_sap3/_1623_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__3182_ heichips25_sap3/_0791_ heichips25_sap3/_0792_ heichips25_sap3/_0790_
+ heichips25_sap3/_0795_ VPWR VGND heichips25_sap3/_0793_ sg13g2_nand4_1
XFILLER_44_377 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2133_ heichips25_sap3/_1554_ heichips25_sap3__4065_/Q heichips25_sap3/_1459_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__2064_ heichips25_sap3/_1468_ heichips25_sap3/_1478_ heichips25_sap3/_1485_
+ VPWR VGND sg13g2_nor2_1
XFILLER_12_230 VPWR VGND sg13g2_decap_4
XFILLER_8_201 VPWR VGND sg13g2_fill_2
XFILLER_9_713 VPWR VGND sg13g2_fill_2
XFILLER_9_735 VPWR VGND sg13g2_decap_4
XFILLER_8_223 VPWR VGND sg13g2_fill_2
XFILLER_12_285 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2966_ heichips25_sap3/net70 heichips25_sap3/net275 heichips25_sap3/_0603_
+ heichips25_sap3/_0047_ VPWR VGND sg13g2_a21o_1
XFILLER_5_996 VPWR VGND sg13g2_decap_8
XFILLER_5_78 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2897_ heichips25_sap3/net69 heichips25_sap3/net281 heichips25_sap3/_0537_
+ heichips25_sap3/_0044_ VPWR VGND sg13g2_a21o_1
Xheichips25_can_lehmann_fsm__2792__623 VPWR VGND net622 sg13g2_tiehi
XFILLER_39_116 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3518_ heichips25_sap3/_0967_ heichips25_sap3/_0970_ heichips25_sap3/net96
+ heichips25_sap3/_1111_ VPWR VGND sg13g2_nand3_1
XFILLER_47_160 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3449_ heichips25_sap3/_1054_ heichips25_sap3/net122 heichips25_sap3/net62
+ VPWR VGND sg13g2_nand2_1
XFILLER_39_1017 VPWR VGND sg13g2_fill_1
XFILLER_36_856 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2670_ heichips25_can_lehmann_fsm/net484 VPWR heichips25_can_lehmann_fsm/_0801_
+ VGND heichips25_can_lehmann_fsm/net915 heichips25_can_lehmann_fsm/net420 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__1621_ VPWR heichips25_can_lehmann_fsm/_0945_ heichips25_can_lehmann_fsm/net879
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__1552_ VPWR heichips25_can_lehmann_fsm/_0876_ heichips25_can_lehmann_fsm/net1129
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__2838__531 VPWR VGND net530 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2104_ heichips25_can_lehmann_fsm/_0444_ heichips25_can_lehmann_fsm/net187
+ heichips25_can_lehmann_fsm/_0443_ heichips25_can_lehmann_fsm/_0304_ heichips25_can_lehmann_fsm/net1262
+ VPWR VGND sg13g2_a22oi_1
XFILLER_49_18 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2035_ heichips25_can_lehmann_fsm/_0385_ heichips25_can_lehmann_fsm/net185
+ heichips25_can_lehmann_fsm/_0384_ VPWR VGND sg13g2_nand2_1
Xheichips25_can_lehmann_fsm__2937_ net587 VGND VPWR heichips25_can_lehmann_fsm/_0162_
+ heichips25_can_lehmann_fsm__2937_/Q clknet_leaf_17_clk sg13g2_dfrbpq_1
XFILLER_38_193 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2868_ net759 VGND VPWR heichips25_can_lehmann_fsm/_0093_
+ heichips25_can_lehmann_fsm__2868_/Q clknet_leaf_20_clk sg13g2_dfrbpq_1
XFILLER_41_303 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1819_ heichips25_can_lehmann_fsm/_0986_ heichips25_can_lehmann_fsm/_0988_
+ heichips25_can_lehmann_fsm/_1122_ heichips25_can_lehmann_fsm/_1135_ VPWR VGND sg13g2_mux2_1
Xheichips25_can_lehmann_fsm__2799_ net608 VGND VPWR heichips25_can_lehmann_fsm/net1265
+ heichips25_can_lehmann_fsm__2799_/Q clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_14_76 VPWR VGND sg13g2_fill_2
XFILLER_6_727 VPWR VGND sg13g2_fill_1
XFILLER_5_226 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2820_ VGND VPWR heichips25_sap3/net289 heichips25_sap3/_0462_ heichips25_sap3/_0464_
+ heichips25_sap3/_0463_ sg13g2_a21oi_1
Xheichips25_sap3__2751_ heichips25_sap3/_0386_ VPWR heichips25_sap3/_0397_ VGND heichips25_sap3/_0385_
+ heichips25_sap3/_0396_ sg13g2_o21ai_1
XFILLER_30_86 VPWR VGND sg13g2_decap_8
XFILLER_2_944 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2682_ heichips25_sap3/_0331_ VPWR heichips25_sap3/_0027_ VGND heichips25_sap3/_1383_
+ heichips25_sap3/net213 sg13g2_o21ai_1
XFILLER_18_801 VPWR VGND sg13g2_fill_1
XFILLER_17_311 VPWR VGND sg13g2_decap_4
XFILLER_18_823 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3303_ heichips25_sap3/_0854_ VPWR heichips25_sap3/_0914_ VGND heichips25_sap3/_0841_
+ heichips25_sap3/_0902_ sg13g2_o21ai_1
XFILLER_17_344 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3234_ heichips25_sap3/_0718_ heichips25_sap3/_0762_ heichips25_sap3__3948_/Q
+ heichips25_sap3/_0847_ VPWR VGND sg13g2_nand3_1
XFILLER_44_163 VPWR VGND sg13g2_fill_1
XFILLER_44_152 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3165_ heichips25_sap3/_0778_ heichips25_sap3/_0775_ heichips25_sap3/_0776_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__2116_ heichips25_sap3/_1537_ heichips25_sap3/_1513_ heichips25_sap3/_1532_
+ VPWR VGND sg13g2_nand2_1
XFILLER_33_859 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3096_ heichips25_sap3/net222 heichips25_sap3/_0708_ heichips25_sap3/_0709_
+ VPWR VGND sg13g2_nor2_1
XFILLER_9_521 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2047_ heichips25_sap3/net252 heichips25_sap3/net253 heichips25_sap3/_1468_
+ VPWR VGND sg13g2_xor2_1
XFILLER_9_576 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3998_ heichips25_sap3/net439 VGND VPWR heichips25_sap3/_0139_ heichips25_sap3__3998_/Q
+ clkload18/A sg13g2_dfrbpq_1
Xheichips25_sap3__2949_ heichips25_sap3/_0587_ heichips25_sap3/_0585_ heichips25_sap3/_0586_
+ VPWR VGND sg13g2_xnor2_1
Xheichips25_can_lehmann_fsm__2722_ heichips25_can_lehmann_fsm/net478 VPWR heichips25_can_lehmann_fsm/_0827_
+ VGND heichips25_can_lehmann_fsm/net1172 heichips25_can_lehmann_fsm/net369 sg13g2_o21ai_1
XFILLER_24_826 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2653_ VGND VPWR heichips25_can_lehmann_fsm/_0882_ heichips25_can_lehmann_fsm/net381
+ heichips25_can_lehmann_fsm/_0226_ heichips25_can_lehmann_fsm/_0792_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__1604_ VPWR heichips25_can_lehmann_fsm/_0928_ heichips25_can_lehmann_fsm/net1049
+ VGND sg13g2_inv_1
XFILLER_24_848 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2584_ heichips25_can_lehmann_fsm/net476 VPWR heichips25_can_lehmann_fsm/_0758_
+ VGND heichips25_can_lehmann_fsm__2966_/Q heichips25_can_lehmann_fsm/net358 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2961__781 VPWR VGND net780 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__1535_ VPWR heichips25_can_lehmann_fsm/_0859_ heichips25_can_lehmann_fsm/net1151
+ VGND sg13g2_inv_1
XFILLER_31_391 VPWR VGND sg13g2_fill_2
XFILLER_2_207 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2018_ heichips25_can_lehmann_fsm/_0371_ heichips25_can_lehmann_fsm/net184
+ heichips25_can_lehmann_fsm/_0370_ heichips25_can_lehmann_fsm/net191 heichips25_can_lehmann_fsm/net1249
+ VPWR VGND sg13g2_a22oi_1
XFILLER_27_631 VPWR VGND sg13g2_fill_1
XFILLER_27_675 VPWR VGND sg13g2_fill_1
XFILLER_26_185 VPWR VGND sg13g2_fill_1
XFILLER_42_667 VPWR VGND sg13g2_fill_1
XFILLER_41_41 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3921_ heichips25_sap3/net450 VGND VPWR heichips25_sap3/_0062_ heichips25_sap3__3921_/Q
+ heichips25_sap3__3921_/CLK sg13g2_dfrbpq_1
XFILLER_6_524 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3852_ heichips25_sap3/_1349_ VPWR heichips25_sap3/_1352_ VGND heichips25_sap3__4047_/Q
+ heichips25_sap3/_1351_ sg13g2_o21ai_1
Xheichips25_sap3__2803_ heichips25_sap3/_0372_ heichips25_sap3/net254 heichips25_sap3/_0448_
+ VPWR VGND sg13g2_xor2_1
Xheichips25_sap3__3783_ VPWR VGND heichips25_sap3/_1293_ heichips25_sap3/net339 heichips25_sap3/_1287_
+ heichips25_sap3/_1385_ heichips25_sap3/_1294_ heichips25_sap3/net290 sg13g2_a221oi_1
XFILLER_2_730 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2734_ heichips25_sap3/_0351_ heichips25_sap3/_0353_ heichips25_sap3/_0380_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__2665_ VPWR VGND heichips25_sap3/_1907_ heichips25_sap3/net67 heichips25_sap3/_1904_
+ heichips25_sap3/_1385_ uio_oe_sap3\[1\] heichips25_sap3/net89 sg13g2_a221oi_1
Xheichips25_sap3__2596_ heichips25_sap3/_0257_ heichips25_sap3/_0258_ heichips25_sap3/_0261_
+ heichips25_sap3/_0268_ uio_out_sap3\[2\] VPWR VGND sg13g2_or4_1
Xheichips25_sap3__3217_ heichips25_sap3/_0826_ heichips25_sap3/_0827_ heichips25_sap3/_0825_
+ heichips25_sap3/_0830_ VPWR VGND heichips25_sap3/_0828_ sg13g2_nand4_1
XFILLER_20_306 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3148_ heichips25_sap3/_0761_ heichips25_sap3/net145 heichips25_sap3__3955_/Q
+ heichips25_sap3/net108 heichips25_sap3__3947_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_32_144 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3079_ heichips25_sap3/_1697_ heichips25_sap3/_0648_ heichips25_sap3/_0683_
+ heichips25_sap3/_0687_ heichips25_sap3/_0692_ VPWR VGND sg13g2_or4_1
XFILLER_13_391 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_fanout405 heichips25_can_lehmann_fsm/net407 heichips25_can_lehmann_fsm/net405
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout427 heichips25_can_lehmann_fsm/net429 heichips25_can_lehmann_fsm/net427
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout416 heichips25_can_lehmann_fsm/net420 heichips25_can_lehmann_fsm/net416
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm__2705_ VGND VPWR heichips25_can_lehmann_fsm/_0869_ heichips25_can_lehmann_fsm/net428
+ heichips25_can_lehmann_fsm/_0252_ heichips25_can_lehmann_fsm/_0818_ sg13g2_a21oi_1
XFILLER_24_612 VPWR VGND sg13g2_fill_2
XFILLER_23_100 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2636_ heichips25_can_lehmann_fsm/net465 VPWR heichips25_can_lehmann_fsm/_0784_
+ VGND heichips25_can_lehmann_fsm/net964 heichips25_can_lehmann_fsm/net357 sg13g2_o21ai_1
XFILLER_24_678 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2567_ VGND VPWR heichips25_can_lehmann_fsm/_0906_ heichips25_can_lehmann_fsm/net418
+ heichips25_can_lehmann_fsm/_0183_ heichips25_can_lehmann_fsm/_0749_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2498_ heichips25_can_lehmann_fsm/net467 VPWR heichips25_can_lehmann_fsm/_0715_
+ VGND heichips25_can_lehmann_fsm__2924_/Q heichips25_can_lehmann_fsm/net391 sg13g2_o21ai_1
Xheichips25_sap3__2450_ heichips25_sap3/_1856_ heichips25_sap3/_1864_ uio_out_sap3\[4\]
+ VPWR VGND heichips25_sap3/_1852_ sg13g2_nand3b_1
Xheichips25_sap3__2381_ heichips25_sap3/_1442_ heichips25_sap3/_1495_ heichips25_sap3/net226
+ heichips25_sap3/_1801_ VPWR VGND sg13g2_nor3_1
XFILLER_36_63 VPWR VGND sg13g2_decap_4
XFILLER_43_943 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__4051_ heichips25_sap3/net451 VGND VPWR heichips25_sap3/_0192_ heichips25_sap3__4051_/Q
+ clknet_leaf_23_clk sg13g2_dfrbpq_1
XFILLER_14_100 VPWR VGND sg13g2_decap_8
XFILLER_14_122 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3002_ heichips25_sap3__3918_/Q heichips25_sap3/net201 heichips25_sap3/_0628_
+ VPWR VGND sg13g2_nor2_1
XFILLER_30_659 VPWR VGND sg13g2_decap_8
Xinput16 uio_in[5] net16 VPWR VGND sg13g2_buf_1
XFILLER_6_310 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3904_ heichips25_sap3/net455 VGND VPWR heichips25_sap3/_0045_ heichips25_sap3__3904_/Q
+ clkload26/A sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2975__725 VPWR VGND net724 sg13g2_tiehi
Xheichips25_sap3__3835_ heichips25_sap3/_1337_ heichips25_sap3/_1338_ heichips25_sap3/_1336_
+ heichips25_sap3/_1340_ VPWR VGND heichips25_sap3/_1339_ sg13g2_nand4_1
XFILLER_7_899 VPWR VGND sg13g2_decap_8
XFILLER_7_888 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3766_ heichips25_sap3/_1264_ heichips25_sap3/_1271_ heichips25_sap3/_1278_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__3697_ heichips25_sap3/_1230_ VPWR heichips25_sap3/_0151_ VGND heichips25_sap3/_0755_
+ heichips25_sap3/_1177_ sg13g2_o21ai_1
Xheichips25_sap3__2717_ heichips25_sap3__3916_/Q heichips25_sap3/net286 heichips25_sap3/_0363_
+ VPWR VGND sg13g2_xor2_1
Xheichips25_sap3__2648_ heichips25_sap3/_1618_ heichips25_sap3/_1643_ heichips25_sap3/net237
+ heichips25_sap3/_0315_ VPWR VGND sg13g2_nand3_1
XFILLER_37_247 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2579_ heichips25_sap3/_0248_ heichips25_sap3/_0249_ heichips25_sap3/_0250_
+ heichips25_sap3/_0251_ heichips25_sap3/_0252_ VPWR VGND sg13g2_and4_1
XFILLER_18_461 VPWR VGND sg13g2_decap_8
XFILLER_45_291 VPWR VGND sg13g2_fill_1
XFILLER_33_431 VPWR VGND sg13g2_fill_1
XFILLER_21_626 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2421_ VGND VPWR heichips25_can_lehmann_fsm/_0944_ heichips25_can_lehmann_fsm/net427
+ heichips25_can_lehmann_fsm/_0110_ heichips25_can_lehmann_fsm/_0676_ sg13g2_a21oi_1
XFILLER_20_147 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2352_ heichips25_can_lehmann_fsm/net494 VPWR heichips25_can_lehmann_fsm/_0642_
+ VGND heichips25_can_lehmann_fsm/net857 heichips25_can_lehmann_fsm/net383 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2283_ VGND VPWR heichips25_can_lehmann_fsm/net942 heichips25_can_lehmann_fsm/net171
+ heichips25_can_lehmann_fsm/_0597_ heichips25_can_lehmann_fsm/_0596_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2954__809 VPWR VGND net808 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__1998_ VPWR VGND heichips25_can_lehmann_fsm__2786_/Q heichips25_can_lehmann_fsm/net193
+ heichips25_can_lehmann_fsm/net189 heichips25_can_lehmann_fsm__2784_/Q heichips25_can_lehmann_fsm/_0354_
+ heichips25_can_lehmann_fsm/net198 sg13g2_a221oi_1
XFILLER_37_781 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2619_ VGND VPWR heichips25_can_lehmann_fsm/_0893_ heichips25_can_lehmann_fsm/net417
+ heichips25_can_lehmann_fsm/_0209_ heichips25_can_lehmann_fsm/_0775_ sg13g2_a21oi_1
XFILLER_22_76 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__1950_ VPWR heichips25_sap3/_1376_ heichips25_sap3__4013_/Q VGND
+ sg13g2_inv_1
XFILLER_4_847 VPWR VGND sg13g2_decap_8
XFILLER_3_357 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3620_ heichips25_sap3/net102 heichips25_sap3/_1067_ heichips25_sap3/_1182_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__3551_ heichips25_sap3__3958_/Q heichips25_sap3/_1068_ heichips25_sap3/_1134_
+ heichips25_sap3/_0099_ VPWR VGND sg13g2_mux2_1
Xheichips25_sap3__2502_ heichips25_sap3/_1915_ heichips25_sap3/net76 heichips25_sap3__3988_/Q
+ heichips25_sap3/net83 heichips25_sap3__3964_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3482_ heichips25_sap3/_0086_ heichips25_sap3/_1077_ heichips25_sap3/_1080_
+ heichips25_sap3/net57 heichips25_sap3/_1419_ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2433_ heichips25_sap3/_1845_ heichips25_sap3/_1847_ heichips25_sap3/_1848_
+ VPWR VGND sg13g2_and2_1
XFILLER_35_707 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2364_ VGND VPWR heichips25_sap3/_1449_ heichips25_sap3/_1782_ heichips25_sap3/_1785_
+ heichips25_sap3/_1784_ sg13g2_a21oi_1
Xheichips25_sap3__2295_ heichips25_sap3/_1491_ heichips25_sap3/_1538_ heichips25_sap3/net256
+ heichips25_sap3/_1716_ VPWR VGND heichips25_sap3/_1568_ sg13g2_nand4_1
Xheichips25_sap3__4034_ heichips25_sap3/net458 VGND VPWR heichips25_sap3/_0175_ heichips25_sap3__4034_/Q
+ clknet_leaf_1_clk sg13g2_dfrbpq_1
XFILLER_42_250 VPWR VGND sg13g2_decap_8
Xclkbuf_4_15_0_heichips25_sap3\_sap_3_inst.alu_inst.clk clknet_0_heichips25_sap3\/sap_3_inst.alu_inst.clk
+ clknet_4_15_0_heichips25_sap3\/sap_3_inst.alu_inst.clk VPWR VGND sg13g2_buf_8
Xheichips25_can_lehmann_fsm_hold880 heichips25_can_lehmann_fsm__2882_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net879 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold891 heichips25_can_lehmann_fsm/_0212_ VPWR VGND heichips25_can_lehmann_fsm/net890
+ sg13g2_dlygate4sd3_1
XFILLER_11_670 VPWR VGND sg13g2_decap_4
XFILLER_10_191 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__3036__534 VPWR VGND net533 sg13g2_tiehi
Xheichips25_sap3__3818_ VPWR VGND heichips25_sap3__4024_/Q heichips25_sap3/_1324_
+ heichips25_sap3/_1270_ heichips25_sap3__3984_/Q heichips25_sap3/_1325_ heichips25_sap3/_1259_
+ sg13g2_a221oi_1
Xheichips25_sap3__3749_ heichips25_sap3/_1257_ heichips25_sap3/_1260_ heichips25_sap3/_1261_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_can_lehmann_fsm__2970_ net744 VGND VPWR heichips25_can_lehmann_fsm/net888
+ heichips25_can_lehmann_fsm__2970_/Q clknet_leaf_20_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1921_ VGND VPWR heichips25_can_lehmann_fsm/_1223_ heichips25_can_lehmann_fsm/_1224_
+ heichips25_can_lehmann_fsm/_1234_ heichips25_can_lehmann_fsm/_1233_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__1852_ heichips25_can_lehmann_fsm/_1168_ heichips25_can_lehmann_fsm/net297
+ heichips25_can_lehmann_fsm__2890_/Q heichips25_can_lehmann_fsm/net307 heichips25_can_lehmann_fsm__2938_/Q
+ VPWR VGND sg13g2_a22oi_1
X_17_ net518 uio_out_sap3\[3\] net504 net30 VPWR VGND sg13g2_mux2_1
Xheichips25_can_lehmann_fsm__1783_ heichips25_can_lehmann_fsm__2807_/Q heichips25_can_lehmann_fsm__2806_/Q
+ heichips25_can_lehmann_fsm/_1098_ heichips25_can_lehmann_fsm/_1099_ VPWR VGND sg13g2_nor3_1
Xheichips25_sap3_rebuffer829 net829 heichips25_sap3/net828 VPWR VGND sg13g2_buf_1
Xheichips25_sap3_fanout106 heichips25_sap3/_0758_ heichips25_sap3/net106 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout128 heichips25_sap3/net130 heichips25_sap3/net128 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout117 heichips25_sap3/net118 heichips25_sap3/net117 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout139 heichips25_sap3/_0768_ heichips25_sap3/net139 VPWR VGND
+ sg13g2_buf_1
Xheichips25_can_lehmann_fsm_hold1218 heichips25_can_lehmann_fsm__2815_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1217 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1207 heichips25_can_lehmann_fsm/_0042_ VPWR VGND heichips25_can_lehmann_fsm/net1206
+ sg13g2_dlygate4sd3_1
XFILLER_34_795 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_hold1229 heichips25_can_lehmann_fsm/_0017_ VPWR VGND heichips25_can_lehmann_fsm/net1228
+ sg13g2_dlygate4sd3_1
Xheichips25_sap3_hold927 heichips25_sap3/_0176_ VPWR VGND heichips25_sap3/net926 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__2404_ heichips25_can_lehmann_fsm/net473 VPWR heichips25_can_lehmann_fsm/_0668_
+ VGND heichips25_can_lehmann_fsm/net1126 heichips25_can_lehmann_fsm/net401 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2335_ VGND VPWR heichips25_can_lehmann_fsm/_0968_ heichips25_can_lehmann_fsm/net408
+ heichips25_can_lehmann_fsm/_0067_ heichips25_can_lehmann_fsm/_0633_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2266_ heichips25_can_lehmann_fsm/_0583_ heichips25_can_lehmann_fsm/net1194
+ heichips25_can_lehmann_fsm/_1045_ VPWR VGND sg13g2_xnor2_1
Xheichips25_can_lehmann_fsm__2197_ heichips25_can_lehmann_fsm/_0529_ heichips25_can_lehmann_fsm/net164
+ heichips25_can_lehmann_fsm/_0528_ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__2080_ heichips25_sap3/_1501_ heichips25_sap3/net272 heichips25_sap3/net269
+ VPWR VGND sg13g2_nand2_1
XFILLER_12_412 VPWR VGND sg13g2_decap_8
XFILLER_25_773 VPWR VGND sg13g2_fill_2
XFILLER_8_416 VPWR VGND sg13g2_decap_8
XFILLER_12_489 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2779__649 VPWR VGND net648 sg13g2_tiehi
Xheichips25_sap3__2982_ heichips25_sap3/_0051_ heichips25_sap3/_0614_ heichips25_sap3/_0615_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__1933_ VPWR heichips25_sap3/_1359_ heichips25_sap3/net1064 VGND sg13g2_inv_1
XFILLER_4_655 VPWR VGND sg13g2_fill_2
XFILLER_3_154 VPWR VGND sg13g2_decap_8
XFILLER_3_132 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3603_ heichips25_sap3/_1175_ heichips25_sap3/_1063_ heichips25_sap3/_1174_
+ VPWR VGND sg13g2_nand2_1
XFILLER_0_850 VPWR VGND sg13g2_fill_2
XFILLER_39_309 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3534_ net43 uio_oe_sap3\[6\] heichips25_sap3/_1087_ heichips25_sap3/_1125_
+ VPWR VGND sg13g2_mux2_1
Xheichips25_sap3__3465_ heichips25_sap3/net45 VPWR heichips25_sap3/_1067_ VGND heichips25_sap3/net119
+ heichips25_sap3/_0957_ sg13g2_o21ai_1
XFILLER_47_342 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2416_ heichips25_sap3/_1833_ heichips25_sap3/net155 heichips25_sap3/_1832_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__3396_ heichips25_sap3/net121 VPWR heichips25_sap3/_1004_ VGND heichips25_sap3/net126
+ heichips25_sap3/_1003_ sg13g2_o21ai_1
Xheichips25_sap3__2347_ heichips25_sap3/_1766_ heichips25_sap3/_1767_ heichips25_sap3/_1452_
+ heichips25_sap3/_1768_ VPWR VGND sg13g2_nand3_1
Xheichips25_sap3__2278_ VPWR VGND heichips25_sap3/net262 heichips25_sap3/_1574_ heichips25_sap3/_1662_
+ heichips25_sap3/_1537_ heichips25_sap3/_1699_ heichips25_sap3/_1555_ sg13g2_a221oi_1
XFILLER_31_710 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__4017_ heichips25_sap3/net440 VGND VPWR heichips25_sap3/_0158_ heichips25_sap3__4017_/Q
+ heichips25_sap3__4017_/CLK sg13g2_dfrbpq_1
XFILLER_15_272 VPWR VGND sg13g2_fill_2
XFILLER_31_732 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2120_ heichips25_can_lehmann_fsm/_0458_ VPWR heichips25_can_lehmann_fsm/_0459_
+ VGND heichips25_can_lehmann_fsm__2879_/Q heichips25_can_lehmann_fsm/net335 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2051_ heichips25_can_lehmann_fsm/_0399_ heichips25_can_lehmann_fsm__2797_/Q
+ heichips25_can_lehmann_fsm/net346 VPWR VGND sg13g2_xnor2_1
Xheichips25_can_lehmann_fsm__2953_ net812 VGND VPWR heichips25_can_lehmann_fsm/_0178_
+ heichips25_can_lehmann_fsm__2953_/Q clknet_leaf_9_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1904_ heichips25_can_lehmann_fsm/_1217_ heichips25_can_lehmann_fsm__3009_/Q
+ heichips25_can_lehmann_fsm/net318 VPWR VGND sg13g2_nand2_1
Xheichips25_can_lehmann_fsm__2884_ net727 VGND VPWR heichips25_can_lehmann_fsm/_0109_
+ heichips25_can_lehmann_fsm__2884_/Q clknet_leaf_11_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1835_ VGND VPWR heichips25_can_lehmann_fsm/_1054_ heichips25_can_lehmann_fsm/_1140_
+ heichips25_can_lehmann_fsm/_1151_ heichips25_can_lehmann_fsm/_1150_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm_hold1004 heichips25_can_lehmann_fsm__2887_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1003 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__1766_ heichips25_can_lehmann_fsm/_1083_ heichips25_can_lehmann_fsm/_1032_
+ heichips25_can_lehmann_fsm__2801_/Q heichips25_can_lehmann_fsm/_1031_ heichips25_can_lehmann_fsm/net350
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm_hold1026 heichips25_can_lehmann_fsm__2943_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1025 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1015 heichips25_can_lehmann_fsm/_0163_ VPWR VGND heichips25_can_lehmann_fsm/net1014
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__1697_ heichips25_can_lehmann_fsm/_1018_ heichips25_can_lehmann_fsm/_1019_
+ heichips25_can_lehmann_fsm/_1017_ heichips25_can_lehmann_fsm/_1021_ VPWR VGND heichips25_can_lehmann_fsm/_1020_
+ sg13g2_nand4_1
Xheichips25_can_lehmann_fsm_hold1037 heichips25_can_lehmann_fsm/_0182_ VPWR VGND heichips25_can_lehmann_fsm/net1036
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1048 heichips25_can_lehmann_fsm__2925_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1047 sg13g2_dlygate4sd3_1
XFILLER_10_905 VPWR VGND sg13g2_fill_1
XFILLER_21_297 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2318_ heichips25_can_lehmann_fsm/net473 VPWR heichips25_can_lehmann_fsm/_0625_
+ VGND heichips25_can_lehmann_fsm/net1204 heichips25_can_lehmann_fsm/net401 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2249_ VGND VPWR heichips25_can_lehmann_fsm/net210 heichips25_can_lehmann_fsm/_0568_
+ heichips25_can_lehmann_fsm/_0045_ heichips25_can_lehmann_fsm/_0569_ sg13g2_a21oi_1
XFILLER_0_135 VPWR VGND sg13g2_decap_8
XFILLER_1_636 VPWR VGND sg13g2_fill_1
XFILLER_1_669 VPWR VGND sg13g2_fill_2
XFILLER_0_146 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3250_ VGND VPWR heichips25_sap3/_0863_ heichips25_sap3/net166 heichips25_sap3/_0731_
+ sg13g2_or2_1
XFILLER_28_53 VPWR VGND sg13g2_fill_2
XFILLER_45_846 VPWR VGND sg13g2_fill_2
XFILLER_44_312 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2201_ VGND VPWR heichips25_sap3/_1622_ heichips25_sap3/_1620_ heichips25_sap3/_1618_
+ sg13g2_or2_1
XFILLER_17_526 VPWR VGND sg13g2_decap_8
XFILLER_29_386 VPWR VGND sg13g2_fill_2
XFILLER_45_879 VPWR VGND sg13g2_fill_1
XFILLER_45_857 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3181_ heichips25_sap3/_0790_ heichips25_sap3/_0791_ heichips25_sap3/_0792_
+ heichips25_sap3/_0793_ heichips25_sap3/_0794_ VPWR VGND sg13g2_and4_1
Xheichips25_sap3__2132_ heichips25_sap3/_1553_ heichips25_sap3/_1551_ heichips25_sap3/_1463_
+ heichips25_sap3/_1546_ heichips25_sap3/net246 VPWR VGND sg13g2_a22oi_1
XFILLER_25_570 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2063_ heichips25_sap3/_1473_ heichips25_sap3/_1482_ heichips25_sap3/_1483_
+ heichips25_sap3/_1484_ VPWR VGND sg13g2_nor3_1
XFILLER_9_758 VPWR VGND sg13g2_fill_2
XFILLER_8_279 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2965_ heichips25_sap3/_0440_ heichips25_sap3/_0584_ heichips25_sap3/_0602_
+ heichips25_sap3/_0603_ VPWR VGND sg13g2_nor3_1
XFILLER_4_452 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2896_ heichips25_sap3/net69 heichips25_sap3/_0518_ heichips25_sap3/_0536_
+ heichips25_sap3/_0537_ VPWR VGND sg13g2_nor3_1
Xheichips25_sap3__3517_ heichips25_sap3__3951_/Q heichips25_sap3/net109 heichips25_sap3/_1110_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__3448_ heichips25_sap3/net119 heichips25_sap3/net59 heichips25_sap3/_1053_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__3379_ heichips25_sap3/_0987_ heichips25_sap3/net139 heichips25_sap3__3976_/Q
+ heichips25_sap3/net143 heichips25_sap3__3984_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_35_334 VPWR VGND sg13g2_decap_8
XFILLER_35_367 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1620_ VPWR heichips25_can_lehmann_fsm/_0944_ heichips25_can_lehmann_fsm/net976
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__1551_ VPWR heichips25_can_lehmann_fsm/_0875_ heichips25_can_lehmann_fsm/net853
+ VGND sg13g2_inv_1
Xclkbuf_5_11__f_heichips25_sap3\_sap_3_inst.alu_inst.clk clkload20/A clknet_4_5_0_heichips25_sap3\/sap_3_inst.alu_inst.clk
+ VPWR VGND sg13g2_buf_16
Xheichips25_can_lehmann_fsm__2103_ heichips25_can_lehmann_fsm/_0443_ heichips25_can_lehmann_fsm/_0442_
+ heichips25_can_lehmann_fsm/_1060_ VPWR VGND sg13g2_nand2b_1
XFILLER_7_290 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2034_ heichips25_can_lehmann_fsm/_0384_ heichips25_can_lehmann_fsm/_0979_
+ heichips25_can_lehmann_fsm/_1073_ VPWR VGND sg13g2_xnor2_1
XFILLER_38_172 VPWR VGND sg13g2_decap_8
XFILLER_38_161 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2936_ net591 VGND VPWR heichips25_can_lehmann_fsm/_0161_
+ heichips25_can_lehmann_fsm__2936_/Q clknet_leaf_17_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2867_ net761 VGND VPWR heichips25_can_lehmann_fsm/_0092_
+ heichips25_can_lehmann_fsm__2867_/Q clknet_leaf_14_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2798_ net610 VGND VPWR heichips25_can_lehmann_fsm/net1267
+ heichips25_can_lehmann_fsm__2798_/Q clknet_leaf_3_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1818_ heichips25_can_lehmann_fsm/_1114_ heichips25_can_lehmann_fsm/_1122_
+ heichips25_can_lehmann_fsm/_1134_ VPWR VGND sg13g2_nor2b_1
XFILLER_41_348 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1749_ VGND VPWR heichips25_can_lehmann_fsm/_1069_ heichips25_can_lehmann_fsm__2786_/Q
+ heichips25_can_lehmann_fsm__2787_/Q sg13g2_or2_1
XFILLER_14_33 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2750_ VGND VPWR heichips25_sap3/_0355_ heichips25_sap3/_0394_ heichips25_sap3/_0396_
+ heichips25_sap3/_0395_ sg13g2_a21oi_1
Xheichips25_sap3__2681_ heichips25_sap3/_0331_ heichips25_sap3__3886_/Q heichips25_sap3/net213
+ VPWR VGND sg13g2_nand2_1
XFILLER_39_85 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3302_ heichips25_sap3/_0891_ VPWR heichips25_sap3/_0073_ VGND heichips25_sap3/_0908_
+ heichips25_sap3/_0913_ sg13g2_o21ai_1
XFILLER_18_813 VPWR VGND sg13g2_fill_2
XFILLER_44_120 VPWR VGND sg13g2_fill_2
XFILLER_18_879 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3233_ heichips25_sap3/_0680_ heichips25_sap3/_0718_ heichips25_sap3__3940_/Q
+ heichips25_sap3/_0846_ VPWR VGND sg13g2_nand3_1
XFILLER_45_676 VPWR VGND sg13g2_fill_1
XFILLER_17_356 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3164_ heichips25_sap3/_0775_ heichips25_sap3/_0776_ heichips25_sap3/_0777_
+ VPWR VGND sg13g2_and2_1
XFILLER_33_805 VPWR VGND sg13g2_decap_8
XFILLER_33_838 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2115_ heichips25_sap3/net243 heichips25_sap3/_1531_ heichips25_sap3/_1536_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__3095_ heichips25_sap3/_1503_ heichips25_sap3/net242 heichips25_sap3/_0295_
+ heichips25_sap3/_0708_ VPWR VGND sg13g2_nor3_1
XFILLER_13_540 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2046_ heichips25_sap3/net253 heichips25_sap3/net252 heichips25_sap3/_1467_
+ VPWR VGND sg13g2_nor2b_1
Xheichips25_can_lehmann_fsm__2904__688 VPWR VGND net687 sg13g2_tiehi
XFILLER_9_555 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3997_ heichips25_sap3/net438 VGND VPWR heichips25_sap3/_0138_ heichips25_sap3__3997_/Q
+ heichips25_sap3__4014_/CLK sg13g2_dfrbpq_1
Xheichips25_sap3__2948_ heichips25_sap3/_0586_ heichips25_sap3/_1374_ heichips25_sap3/net212
+ VPWR VGND sg13g2_xnor2_1
XFILLER_4_271 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2879_ heichips25_sap3/net159 VPWR heichips25_sap3/_0520_ VGND heichips25_sap3/net281
+ heichips25_sap3__3919_/Q sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2721_ VGND VPWR heichips25_can_lehmann_fsm/_0865_ heichips25_can_lehmann_fsm/net410
+ heichips25_can_lehmann_fsm/_0260_ heichips25_can_lehmann_fsm/_0826_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2652_ heichips25_can_lehmann_fsm/net492 VPWR heichips25_can_lehmann_fsm/_0792_
+ VGND heichips25_can_lehmann_fsm__3000_/Q heichips25_can_lehmann_fsm/net381 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__1603_ VPWR heichips25_can_lehmann_fsm/_0927_ heichips25_can_lehmann_fsm/net861
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__2583_ VGND VPWR heichips25_can_lehmann_fsm/_0902_ heichips25_can_lehmann_fsm/net410
+ heichips25_can_lehmann_fsm/_0191_ heichips25_can_lehmann_fsm/_0757_ sg13g2_a21oi_1
XFILLER_32_860 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1534_ VPWR heichips25_can_lehmann_fsm/_0858_ heichips25_can_lehmann_fsm/net1147
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__2805__597 VPWR VGND net596 sg13g2_tiehi
XFILLER_2_219 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2017_ heichips25_can_lehmann_fsm/_0370_ heichips25_can_lehmann_fsm/net1259
+ heichips25_can_lehmann_fsm/_1070_ VPWR VGND sg13g2_xnor2_1
XFILLER_18_109 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2919_ net657 VGND VPWR heichips25_can_lehmann_fsm/_0144_
+ heichips25_can_lehmann_fsm__2919_/Q clknet_leaf_19_clk sg13g2_dfrbpq_1
XFILLER_15_805 VPWR VGND sg13g2_fill_1
XFILLER_25_54 VPWR VGND sg13g2_decap_8
XFILLER_25_65 VPWR VGND sg13g2_fill_2
XFILLER_10_510 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3920_ heichips25_sap3/net448 VGND VPWR heichips25_sap3/_0061_ heichips25_sap3__3920_/Q
+ heichips25_sap3__3920_/CLK sg13g2_dfrbpq_1
XFILLER_10_565 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3851_ heichips25_sap3/_1350_ VPWR heichips25_sap3/_1351_ VGND heichips25_sap3/net342
+ heichips25_sap3__4054_/Q sg13g2_o21ai_1
Xheichips25_sap3__2802_ VGND VPWR heichips25_sap3/_0447_ heichips25_sap3/_0443_ heichips25_sap3/net288
+ sg13g2_or2_1
Xheichips25_sap3__3782_ VPWR VGND heichips25_sap3__4012_/Q heichips25_sap3/_1292_
+ heichips25_sap3/_1281_ heichips25_sap3__3972_/Q heichips25_sap3/_1293_ heichips25_sap3/_1272_
+ sg13g2_a221oi_1
Xheichips25_sap3__2733_ heichips25_sap3/_0374_ heichips25_sap3/_0375_ heichips25_sap3/_0378_
+ heichips25_sap3/_0379_ VPWR VGND sg13g2_or3_1
XFILLER_29_1028 VPWR VGND sg13g2_fill_1
XFILLER_2_753 VPWR VGND sg13g2_fill_2
XFILLER_2_797 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2664_ VPWR VGND heichips25_sap3/_0198_ heichips25_sap3/net67 heichips25_sap3/_1930_
+ heichips25_sap3/_1392_ uio_oe_sap3\[0\] heichips25_sap3/net92 sg13g2_a221oi_1
XFILLER_49_245 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2595_ VGND VPWR heichips25_sap3/_0264_ heichips25_sap3/_0267_ heichips25_sap3/_0268_
+ heichips25_sap3/net67 sg13g2_a21oi_1
XFILLER_49_289 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3216_ heichips25_sap3/_0825_ heichips25_sap3/_0826_ heichips25_sap3/_0827_
+ heichips25_sap3/_0828_ heichips25_sap3/_0829_ VPWR VGND sg13g2_and4_1
XFILLER_17_186 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3147_ heichips25_sap3/_0697_ heichips25_sap3/_0714_ heichips25_sap3/_0716_
+ heichips25_sap3/_0759_ heichips25_sap3/_0760_ VPWR VGND sg13g2_and4_1
Xheichips25_sap3__3078_ heichips25_sap3/_0686_ heichips25_sap3/_0688_ heichips25_sap3/_0684_
+ heichips25_sap3/_0691_ VPWR VGND sg13g2_nand3_1
Xheichips25_sap3__2029_ heichips25_sap3/_1450_ heichips25_sap3/net260 heichips25_sap3/net259
+ VPWR VGND sg13g2_nand2b_1
XFILLER_12_1021 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm_fanout406 heichips25_can_lehmann_fsm/net407 heichips25_can_lehmann_fsm/net406
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout428 heichips25_can_lehmann_fsm/net429 heichips25_can_lehmann_fsm/net428
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout417 heichips25_can_lehmann_fsm/net419 heichips25_can_lehmann_fsm/net417
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm__2704_ heichips25_can_lehmann_fsm/net497 VPWR heichips25_can_lehmann_fsm/_0818_
+ VGND heichips25_can_lehmann_fsm__3027_/Q heichips25_can_lehmann_fsm/net428 sg13g2_o21ai_1
X_17__519 VPWR VGND net518 sg13g2_tielo
Xheichips25_can_lehmann_fsm__2635_ VGND VPWR heichips25_can_lehmann_fsm/_0889_ heichips25_can_lehmann_fsm/net394
+ heichips25_can_lehmann_fsm/_0217_ heichips25_can_lehmann_fsm/_0783_ sg13g2_a21oi_1
XFILLER_23_145 VPWR VGND sg13g2_fill_2
XFILLER_11_318 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2566_ heichips25_can_lehmann_fsm/net488 VPWR heichips25_can_lehmann_fsm/_0749_
+ VGND heichips25_can_lehmann_fsm/net1109 heichips25_can_lehmann_fsm/net418 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2497_ VGND VPWR heichips25_can_lehmann_fsm/_0923_ heichips25_can_lehmann_fsm/net355
+ heichips25_can_lehmann_fsm/_0148_ heichips25_can_lehmann_fsm/_0714_ sg13g2_a21oi_1
XFILLER_11_78 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2857__782 VPWR VGND net781 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__3049_ net573 VGND VPWR heichips25_can_lehmann_fsm/_0274_
+ heichips25_can_lehmann_fsm__3049_/Q clknet_leaf_13_clk sg13g2_dfrbpq_1
Xheichips25_sap3__2380_ heichips25_sap3/_1752_ heichips25_sap3/_1792_ heichips25_sap3/_1800_
+ uio_out_sap3\[7\] VPWR VGND sg13g2_or3_1
XFILLER_4_1008 VPWR VGND sg13g2_decap_8
XFILLER_28_985 VPWR VGND sg13g2_fill_1
XFILLER_28_974 VPWR VGND sg13g2_decap_8
XFILLER_42_410 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__4050_ heichips25_sap3/net451 VGND VPWR heichips25_sap3/_0191_ heichips25_sap3__4050_/Q
+ clknet_leaf_23_clk sg13g2_dfrbpq_1
XFILLER_43_977 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3001_ heichips25_sap3/_0627_ VPWR heichips25_sap3/_0058_ VGND heichips25_sap3/_1397_
+ heichips25_sap3/net201 sg13g2_o21ai_1
XFILLER_30_638 VPWR VGND sg13g2_decap_8
XFILLER_30_649 VPWR VGND sg13g2_fill_1
Xinput17 uio_in[6] net17 VPWR VGND sg13g2_buf_1
XFILLER_7_823 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3903_ heichips25_sap3/net455 VGND VPWR heichips25_sap3/_0044_ heichips25_sap3__3903_/Q
+ clkload26/A sg13g2_dfrbpq_1
Xheichips25_sap3__3834_ heichips25_sap3/_1339_ heichips25_sap3/_1270_ heichips25_sap3__4026_/Q
+ heichips25_sap3/_1266_ heichips25_sap3__3962_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_6_377 VPWR VGND sg13g2_fill_2
XFILLER_6_366 VPWR VGND sg13g2_fill_2
XFILLER_42_8 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3765_ VGND VPWR heichips25_sap3__3939_/Q heichips25_sap3/_1274_
+ heichips25_sap3/_1277_ heichips25_sap3/net290 sg13g2_a21oi_1
Xheichips25_sap3__3696_ heichips25_sap3/_1230_ heichips25_sap3__4010_/Q heichips25_sap3/_0755_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__2716_ heichips25_sap3/_1381_ heichips25_sap3/_1396_ heichips25_sap3/_0362_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__2647_ heichips25_sap3/_0314_ heichips25_sap3/_1719_ heichips25_sap3/_0312_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_can_lehmann_fsm__2789__629 VPWR VGND net628 sg13g2_tiehi
Xheichips25_sap3__2578_ heichips25_sap3/_1695_ heichips25_sap3/net827 heichips25_sap3__3949_/Q
+ heichips25_sap3/_0251_ VPWR VGND sg13g2_nand3_1
XFILLER_19_941 VPWR VGND sg13g2_decap_8
XFILLER_19_963 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2420_ heichips25_can_lehmann_fsm/net498 VPWR heichips25_can_lehmann_fsm/_0676_
+ VGND heichips25_can_lehmann_fsm/net916 heichips25_can_lehmann_fsm/net427 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2351_ VGND VPWR heichips25_can_lehmann_fsm/_0964_ heichips25_can_lehmann_fsm/net423
+ heichips25_can_lehmann_fsm/_0075_ heichips25_can_lehmann_fsm/_0641_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2282_ VGND VPWR heichips25_can_lehmann_fsm/_1049_ heichips25_can_lehmann_fsm/_0595_
+ heichips25_can_lehmann_fsm/_0596_ heichips25_can_lehmann_fsm/net171 sg13g2_a21oi_1
XFILLER_9_182 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1997_ heichips25_can_lehmann_fsm__2793_/Q heichips25_can_lehmann_fsm/net196
+ heichips25_can_lehmann_fsm/_0353_ VPWR VGND sg13g2_nor2b_1
XFILLER_43_229 VPWR VGND sg13g2_fill_2
XFILLER_25_944 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2618_ heichips25_can_lehmann_fsm/net485 VPWR heichips25_can_lehmann_fsm/_0775_
+ VGND heichips25_can_lehmann_fsm/net984 heichips25_can_lehmann_fsm/net417 sg13g2_o21ai_1
XFILLER_11_126 VPWR VGND sg13g2_fill_2
XFILLER_11_137 VPWR VGND sg13g2_decap_4
XFILLER_11_148 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2549_ VGND VPWR heichips25_can_lehmann_fsm/_0910_ heichips25_can_lehmann_fsm/net364
+ heichips25_can_lehmann_fsm/_0174_ heichips25_can_lehmann_fsm/_0740_ sg13g2_a21oi_1
XFILLER_20_682 VPWR VGND sg13g2_fill_2
XFILLER_22_88 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3550_ heichips25_sap3__3957_/Q heichips25_sap3/_1066_ heichips25_sap3/net56
+ heichips25_sap3/_0098_ VPWR VGND sg13g2_mux2_1
Xheichips25_sap3__3481_ heichips25_sap3/net57 heichips25_sap3/_1079_ heichips25_sap3/_1080_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__2501_ heichips25_sap3/_1914_ heichips25_sap3/net71 heichips25_sap3__3980_/Q
+ heichips25_sap3/net74 heichips25_sap3__4004_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2432_ heichips25_sap3/_1847_ heichips25_sap3/net80 heichips25_sap3__4023_/Q
+ heichips25_sap3/net84 heichips25_sap3__3959_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2363_ heichips25_sap3/_1784_ heichips25_sap3/net220 heichips25_sap3/_1783_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__2294_ heichips25_sap3/_1715_ heichips25_sap3/net248 heichips25_sap3/_1714_
+ VPWR VGND sg13g2_nand2_1
XFILLER_43_741 VPWR VGND sg13g2_fill_2
XFILLER_43_730 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__4033_ heichips25_sap3/net458 VGND VPWR heichips25_sap3/_0174_ heichips25_sap3__4033_/Q
+ clknet_leaf_1_clk sg13g2_dfrbpq_1
XFILLER_42_273 VPWR VGND sg13g2_fill_1
XFILLER_15_487 VPWR VGND sg13g2_decap_8
XFILLER_16_988 VPWR VGND sg13g2_fill_1
XFILLER_8_46 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm_hold870 heichips25_can_lehmann_fsm__2914_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net869 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold881 heichips25_can_lehmann_fsm/_0108_ VPWR VGND heichips25_can_lehmann_fsm/net880
+ sg13g2_dlygate4sd3_1
Xheichips25_sap3__3817_ heichips25_sap3/_1321_ heichips25_sap3/_1322_ heichips25_sap3/_1320_
+ heichips25_sap3/_1324_ VPWR VGND heichips25_sap3/_1323_ sg13g2_nand4_1
Xheichips25_sap3__3748_ heichips25_sap3/_1260_ heichips25_sap3/net1197 heichips25_sap3/net1178
+ VPWR VGND sg13g2_nand2_1
XFILLER_33_4 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3679_ heichips25_sap3/_1221_ heichips25_sap3/net149 uio_oe_sap3\[7\]
+ VPWR VGND sg13g2_nand2b_1
Xheichips25_can_lehmann_fsm__1920_ heichips25_can_lehmann_fsm/_1090_ VPWR heichips25_can_lehmann_fsm/_1233_
+ VGND heichips25_can_lehmann_fsm/net219 heichips25_can_lehmann_fsm/_1232_ sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__1851_ heichips25_can_lehmann_fsm/_1167_ heichips25_can_lehmann_fsm/net311
+ heichips25_can_lehmann_fsm__3010_/Q heichips25_can_lehmann_fsm/net318 heichips25_can_lehmann_fsm__2986_/Q
+ VPWR VGND sg13g2_a22oi_1
X_16_ net517 net44 net504 net29 VPWR VGND sg13g2_mux2_1
Xheichips25_sap3_fanout107 heichips25_sap3/_0758_ heichips25_sap3/net107 VPWR VGND
+ sg13g2_buf_1
Xheichips25_can_lehmann_fsm__1782_ heichips25_can_lehmann_fsm__2805_/Q heichips25_can_lehmann_fsm__2804_/Q
+ heichips25_can_lehmann_fsm__2803_/Q heichips25_can_lehmann_fsm__2802_/Q heichips25_can_lehmann_fsm/_1098_
+ VPWR VGND sg13g2_or4_1
Xheichips25_sap3_fanout118 heichips25_sap3/_0752_ heichips25_sap3/net118 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout129 heichips25_sap3/net130 heichips25_sap3/net129 VPWR VGND
+ sg13g2_buf_1
XFILLER_18_281 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm_hold1219 heichips25_can_lehmann_fsm__2810_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1218 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1208 heichips25_can_lehmann_fsm__2812_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1207 sg13g2_dlygate4sd3_1
XFILLER_33_273 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2403_ VGND VPWR heichips25_can_lehmann_fsm/_0950_ heichips25_can_lehmann_fsm/net364
+ heichips25_can_lehmann_fsm/_0101_ heichips25_can_lehmann_fsm/_0667_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2334_ heichips25_can_lehmann_fsm/net474 VPWR heichips25_can_lehmann_fsm/_0633_
+ VGND heichips25_can_lehmann_fsm/net974 heichips25_can_lehmann_fsm/net403 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2265_ VGND VPWR heichips25_can_lehmann_fsm/net208 heichips25_can_lehmann_fsm/_0581_
+ heichips25_can_lehmann_fsm/_0048_ heichips25_can_lehmann_fsm/_0582_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2196_ heichips25_can_lehmann_fsm/_0528_ heichips25_can_lehmann_fsm/_0974_
+ heichips25_can_lehmann_fsm/_1100_ VPWR VGND sg13g2_xnor2_1
XFILLER_0_339 VPWR VGND sg13g2_decap_8
XFILLER_16_218 VPWR VGND sg13g2_decap_8
XFILLER_17_44 VPWR VGND sg13g2_decap_8
XFILLER_25_741 VPWR VGND sg13g2_fill_1
XFILLER_33_54 VPWR VGND sg13g2_fill_2
XFILLER_33_76 VPWR VGND sg13g2_decap_4
XFILLER_21_991 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2981_ heichips25_sap3/_0615_ heichips25_sap3/net153 heichips25_sap3/_0404_
+ heichips25_sap3/net167 heichips25_sap3/net282 VPWR VGND sg13g2_a22oi_1
XFILLER_3_111 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__1932_ VPWR heichips25_sap3/_1358_ heichips25_sap3__3890_/Q VGND
+ sg13g2_inv_1
XFILLER_4_645 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3602_ heichips25_sap3/_1174_ heichips25_sap3/_0852_ heichips25_sap3/_0888_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__3533_ VGND VPWR heichips25_sap3/net96 heichips25_sap3/_1019_ heichips25_sap3/_1124_
+ heichips25_sap3/_1123_ sg13g2_a21oi_1
XFILLER_3_188 VPWR VGND sg13g2_fill_2
XFILLER_0_840 VPWR VGND sg13g2_fill_1
XFILLER_0_873 VPWR VGND sg13g2_fill_1
XFILLER_48_855 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3464_ heichips25_sap3/_1066_ heichips25_sap3__3941_/Q heichips25_sap3/net58
+ heichips25_sap3/_0082_ VPWR VGND sg13g2_mux2_1
Xheichips25_sap3__3395_ heichips25_sap3/_1003_ heichips25_sap3/_1002_ heichips25_sap3/_0856_
+ VPWR VGND sg13g2_nand2b_1
XFILLER_35_505 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2415_ heichips25_sap3/_1832_ heichips25_sap3__3895_/Q heichips25_sap3/_1788_
+ VPWR VGND sg13g2_nand2_1
XFILLER_35_538 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2346_ heichips25_sap3/_1767_ heichips25_sap3/_1472_ heichips25_sap3/net227
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__2277_ heichips25_sap3/_1697_ VPWR heichips25_sap3/_1698_ VGND heichips25_sap3/net262
+ heichips25_sap3/net230 sg13g2_o21ai_1
Xheichips25_sap3__4016_ heichips25_sap3/net442 VGND VPWR heichips25_sap3/_0157_ heichips25_sap3__4016_/Q
+ heichips25_sap3__4016_/CLK sg13g2_dfrbpq_1
XFILLER_15_295 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_10_clk clknet_2_3__leaf_clk clknet_leaf_10_clk VPWR VGND sg13g2_buf_8
XFILLER_11_490 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2050_ heichips25_can_lehmann_fsm/_0398_ heichips25_can_lehmann_fsm/net186
+ heichips25_can_lehmann_fsm/_0397_ heichips25_can_lehmann_fsm/net190 heichips25_can_lehmann_fsm/net1242
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2914__668 VPWR VGND net667 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2952_ net527 VGND VPWR heichips25_can_lehmann_fsm/_0177_
+ heichips25_can_lehmann_fsm__2952_/Q clknet_leaf_7_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2883_ net729 VGND VPWR heichips25_can_lehmann_fsm/net880
+ heichips25_can_lehmann_fsm__2883_/Q clknet_leaf_11_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1903_ heichips25_can_lehmann_fsm/_1216_ heichips25_can_lehmann_fsm/_0940_
+ heichips25_can_lehmann_fsm/net302 VPWR VGND sg13g2_nand2_1
Xheichips25_can_lehmann_fsm__1834_ VGND VPWR heichips25_can_lehmann_fsm/_1147_ heichips25_can_lehmann_fsm/_1149_
+ heichips25_can_lehmann_fsm/_1150_ heichips25_can_lehmann_fsm/_1143_ sg13g2_a21oi_1
XFILLER_26_527 VPWR VGND sg13g2_decap_4
XFILLER_0_91 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm_hold1005 heichips25_can_lehmann_fsm/_0113_ VPWR VGND heichips25_can_lehmann_fsm/net1004
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__1765_ heichips25_can_lehmann_fsm/_1082_ heichips25_can_lehmann_fsm__2792_/Q
+ heichips25_can_lehmann_fsm/_1037_ VPWR VGND sg13g2_nand2_1
Xheichips25_can_lehmann_fsm_hold1027 heichips25_can_lehmann_fsm/_0168_ VPWR VGND heichips25_can_lehmann_fsm/net1026
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__1696_ VGND VPWR heichips25_can_lehmann_fsm__3016_/Q heichips25_can_lehmann_fsm/net310
+ heichips25_can_lehmann_fsm/_1020_ heichips25_can_lehmann_fsm/net300 sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm_hold1038 heichips25_can_lehmann_fsm__2948_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1037 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1016 heichips25_can_lehmann_fsm__2874_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1015 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1049 heichips25_can_lehmann_fsm/_0151_ VPWR VGND heichips25_can_lehmann_fsm/net1048
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__2317_ heichips25_can_lehmann_fsm/_0624_ net8 net9 VPWR
+ VGND sg13g2_nand2_1
Xheichips25_can_lehmann_fsm__2248_ heichips25_can_lehmann_fsm/net329 VPWR heichips25_can_lehmann_fsm/_0569_
+ VGND heichips25_can_lehmann_fsm/net1195 heichips25_can_lehmann_fsm/net210 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2179_ VGND VPWR heichips25_can_lehmann_fsm/net160 heichips25_can_lehmann_fsm/_0513_
+ heichips25_can_lehmann_fsm/_0030_ heichips25_can_lehmann_fsm/_0514_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2815__577 VPWR VGND net576 sg13g2_tiehi
XFILLER_28_32 VPWR VGND sg13g2_fill_2
XFILLER_29_332 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2200_ heichips25_sap3/_1618_ heichips25_sap3/_1620_ heichips25_sap3/_1621_
+ VPWR VGND sg13g2_nor2_1
XFILLER_17_538 VPWR VGND sg13g2_fill_2
XFILLER_29_365 VPWR VGND sg13g2_decap_8
XFILLER_44_335 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3180_ heichips25_sap3/_0793_ heichips25_sap3/net109 heichips25_sap3__3961_/Q
+ heichips25_sap3/net129 heichips25_sap3__3945_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3_fanout460 heichips25_sap3/net461 heichips25_sap3/net460 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3__2131_ heichips25_sap3/_1552_ heichips25_sap3/net251 heichips25_sap3/net250
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__2062_ heichips25_sap3/_1483_ heichips25_sap3/net258 heichips25_sap3/_1447_
+ heichips25_sap3/net239 VPWR VGND sg13g2_and3_1
XFILLER_25_582 VPWR VGND sg13g2_decap_8
XFILLER_40_541 VPWR VGND sg13g2_fill_1
Xheichips25_sap3_hold1060 heichips25_sap3/_0168_ VPWR VGND heichips25_sap3/net1059
+ sg13g2_dlygate4sd3_1
XFILLER_8_203 VPWR VGND sg13g2_fill_1
XFILLER_9_726 VPWR VGND sg13g2_decap_4
XFILLER_8_225 VPWR VGND sg13g2_fill_1
XFILLER_5_932 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2964_ VPWR VGND heichips25_sap3/_0601_ heichips25_sap3/_0434_ heichips25_sap3/_0600_
+ heichips25_sap3__3914_/Q heichips25_sap3/_0602_ heichips25_sap3/_0436_ sg13g2_a221oi_1
Xheichips25_sap3__2895_ VPWR VGND heichips25_sap3/_0535_ heichips25_sap3/net157 heichips25_sap3/_0534_
+ heichips25_sap3__3911_/Q heichips25_sap3/_0536_ heichips25_sap3/net203 sg13g2_a221oi_1
XFILLER_0_670 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3516_ heichips25_sap3/_0091_ heichips25_sap3/_1107_ heichips25_sap3/_1109_
+ heichips25_sap3/net106 heichips25_sap3/_1373_ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3447_ heichips25_sap3/net105 heichips25_sap3/_0883_ heichips25_sap3/_1052_
+ VPWR VGND sg13g2_nor2_1
XFILLER_36_825 VPWR VGND sg13g2_fill_2
Xclkbuf_4_8_0_heichips25_sap3\_sap_3_inst.alu_inst.clk clknet_0_heichips25_sap3\/sap_3_inst.alu_inst.clk
+ clknet_4_8_0_heichips25_sap3\/sap_3_inst.alu_inst.clk VPWR VGND sg13g2_buf_8
Xheichips25_sap3__3378_ heichips25_sap3/_0986_ heichips25_sap3__3952_/Q heichips25_sap3/net110
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__2329_ heichips25_sap3/_1750_ heichips25_sap3/net71 heichips25_sap3__3978_/Q
+ heichips25_sap3/net216 heichips25_sap3__4010_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_35_379 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1550_ VPWR heichips25_can_lehmann_fsm/_0874_ heichips25_can_lehmann_fsm/net998
+ VGND sg13g2_inv_1
XFILLER_16_571 VPWR VGND sg13g2_decap_8
XFILLER_16_582 VPWR VGND sg13g2_fill_1
XFILLER_31_552 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2102_ heichips25_can_lehmann_fsm__2801_/Q VPWR heichips25_can_lehmann_fsm/_0442_
+ VGND heichips25_can_lehmann_fsm__2800_/Q heichips25_can_lehmann_fsm/_1058_ sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2033_ VPWR VGND heichips25_can_lehmann_fsm/net193 heichips25_can_lehmann_fsm/_0383_
+ heichips25_can_lehmann_fsm/_0382_ heichips25_can_lehmann_fsm/_0379_ heichips25_can_lehmann_fsm/_0015_
+ heichips25_can_lehmann_fsm/_0381_ sg13g2_a221oi_1
Xheichips25_can_lehmann_fsm__2935_ net595 VGND VPWR heichips25_can_lehmann_fsm/net1107
+ heichips25_can_lehmann_fsm__2935_/Q clknet_leaf_16_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2866_ net763 VGND VPWR heichips25_can_lehmann_fsm/_0091_
+ heichips25_can_lehmann_fsm__2866_/Q clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_26_324 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2797_ net612 VGND VPWR heichips25_can_lehmann_fsm/net1220
+ heichips25_can_lehmann_fsm__2797_/Q clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_42_839 VPWR VGND sg13g2_fill_2
XFILLER_14_519 VPWR VGND sg13g2_decap_8
XFILLER_26_379 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1817_ VPWR VGND heichips25_can_lehmann_fsm/_1114_ heichips25_can_lehmann_fsm/_1130_
+ heichips25_can_lehmann_fsm/_1132_ heichips25_can_lehmann_fsm/_1108_ heichips25_can_lehmann_fsm/_1133_
+ heichips25_can_lehmann_fsm/_1123_ sg13g2_a221oi_1
XFILLER_35_891 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1748_ heichips25_can_lehmann_fsm/_1061_ heichips25_can_lehmann_fsm/_1064_
+ heichips25_can_lehmann_fsm/_0981_ heichips25_can_lehmann_fsm/_1068_ VPWR VGND heichips25_can_lehmann_fsm/_1066_
+ sg13g2_nand4_1
XFILLER_14_45 VPWR VGND sg13g2_decap_8
XFILLER_14_78 VPWR VGND sg13g2_fill_1
XFILLER_22_563 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1679_ heichips25_can_lehmann_fsm/_1003_ heichips25_can_lehmann_fsm/net350
+ heichips25_can_lehmann_fsm/net351 heichips25_can_lehmann_fsm/net354 VPWR VGND sg13g2_and3_1
XFILLER_14_89 VPWR VGND sg13g2_fill_2
XFILLER_2_913 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2680_ heichips25_sap3/_0330_ VPWR heichips25_sap3/_0026_ VGND heichips25_sap3/_1367_
+ heichips25_sap3/net213 sg13g2_o21ai_1
XFILLER_2_979 VPWR VGND sg13g2_decap_8
XFILLER_39_75 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3301_ heichips25_sap3/_0913_ heichips25_sap3/_0747_ heichips25_sap3/_0912_
+ VPWR VGND sg13g2_nand2b_1
XFILLER_17_335 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3232_ heichips25_sap3/_0718_ heichips25_sap3/net150 heichips25_sap3__3956_/Q
+ heichips25_sap3/_0845_ VPWR VGND sg13g2_nand3_1
Xheichips25_can_lehmann_fsm__2867__762 VPWR VGND net761 sg13g2_tiehi
Xheichips25_sap3__3163_ heichips25_sap3/_0776_ heichips25_sap3/_1392_ heichips25_sap3/net127
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__2114_ heichips25_sap3/_1535_ heichips25_sap3/_1528_ heichips25_sap3/_1533_
+ VPWR VGND sg13g2_nand2_1
XFILLER_32_338 VPWR VGND sg13g2_decap_4
Xheichips25_sap3_fanout290 heichips25_sap3/_1276_ heichips25_sap3/net290 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3__3094_ heichips25_sap3/_0701_ heichips25_sap3/_0703_ heichips25_sap3/_0704_
+ heichips25_sap3/_0706_ heichips25_sap3/_0707_ VPWR VGND sg13g2_and4_1
XFILLER_9_512 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2045_ heichips25_sap3/_1466_ heichips25_sap3/net247 heichips25_sap3/_1463_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_can_lehmann_fsm__2978__713 VPWR VGND net712 sg13g2_tiehi
XFILLER_40_393 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3996_ heichips25_sap3/net434 VGND VPWR heichips25_sap3/_0137_ heichips25_sap3__3996_/Q
+ heichips25_sap3__3996_/CLK sg13g2_dfrbpq_1
Xheichips25_sap3__2947_ heichips25_sap3/_0575_ VPWR heichips25_sap3/_0585_ VGND heichips25_sap3/_0576_
+ heichips25_sap3/_0578_ sg13g2_o21ai_1
Xheichips25_sap3__2878_ heichips25_sap3/_0519_ heichips25_sap3/_0354_ heichips25_sap3/_0449_
+ VPWR VGND sg13g2_nand2_1
XFILLER_49_983 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2720_ heichips25_can_lehmann_fsm/net478 VPWR heichips25_can_lehmann_fsm/_0826_
+ VGND heichips25_can_lehmann_fsm/net1172 heichips25_can_lehmann_fsm/net410 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2651_ VGND VPWR heichips25_can_lehmann_fsm/_0883_ heichips25_can_lehmann_fsm/net421
+ heichips25_can_lehmann_fsm/_0225_ heichips25_can_lehmann_fsm/_0791_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__1602_ VPWR heichips25_can_lehmann_fsm/_0926_ heichips25_can_lehmann_fsm/net1108
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__2582_ heichips25_can_lehmann_fsm/net476 VPWR heichips25_can_lehmann_fsm/_0757_
+ VGND heichips25_can_lehmann_fsm/net902 heichips25_can_lehmann_fsm/net410 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2799__609 VPWR VGND net608 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__1533_ VPWR heichips25_can_lehmann_fsm/_0857_ heichips25_can_lehmann_fsm/net1117
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__2016_ VPWR VGND heichips25_can_lehmann_fsm/net1246 heichips25_can_lehmann_fsm/net181
+ heichips25_can_lehmann_fsm/net188 heichips25_can_lehmann_fsm/net1240 heichips25_can_lehmann_fsm/_0369_
+ heichips25_can_lehmann_fsm/net197 sg13g2_a221oi_1
Xheichips25_can_lehmann_fsm__2918_ net659 VGND VPWR heichips25_can_lehmann_fsm/_0143_
+ heichips25_can_lehmann_fsm__2918_/Q clknet_leaf_19_clk sg13g2_dfrbpq_1
XFILLER_26_121 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2849_ net797 VGND VPWR heichips25_can_lehmann_fsm/_0074_
+ heichips25_can_lehmann_fsm__2849_/Q clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_26_165 VPWR VGND sg13g2_fill_1
XFILLER_41_179 VPWR VGND sg13g2_decap_4
XFILLER_41_98 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3850_ heichips25_sap3/_1350_ heichips25_sap3/net342 heichips25_sap3__4055_/Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_10_599 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2801_ heichips25_sap3/net154 heichips25_sap3/net64 heichips25_sap3/_0445_
+ heichips25_sap3/_0446_ VPWR VGND sg13g2_or3_1
Xheichips25_sap3__3781_ heichips25_sap3/_1289_ heichips25_sap3/_1290_ heichips25_sap3/_1288_
+ heichips25_sap3/_1292_ VPWR VGND heichips25_sap3/_1291_ sg13g2_nand4_1
Xheichips25_can_lehmann_fsm__3038__791 VPWR VGND net790 sg13g2_tiehi
Xheichips25_sap3__2732_ heichips25_sap3/_0377_ heichips25_sap3/_0366_ heichips25_sap3/_0378_
+ VPWR VGND sg13g2_xor2_1
XFILLER_2_765 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2663_ VGND VPWR heichips25_sap3/_1606_ heichips25_sap3/_0326_ heichips25_sap3/_0006_
+ heichips25_sap3/_0323_ sg13g2_a21oi_1
XFILLER_49_224 VPWR VGND sg13g2_decap_8
XFILLER_2_15 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2594_ heichips25_sap3/_0262_ heichips25_sap3/_0263_ heichips25_sap3/_0265_
+ heichips25_sap3/_0266_ heichips25_sap3/_0267_ VPWR VGND sg13g2_and4_1
XFILLER_49_268 VPWR VGND sg13g2_decap_8
XFILLER_18_600 VPWR VGND sg13g2_fill_1
XFILLER_17_132 VPWR VGND sg13g2_decap_8
XFILLER_17_143 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3215_ heichips25_sap3/_0828_ heichips25_sap3__3963_/Q heichips25_sap3/net145
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__3146_ VPWR VGND heichips25_sap3/_0677_ heichips25_sap3/_0664_ heichips25_sap3/_0676_
+ heichips25_sap3/net241 heichips25_sap3/_0759_ heichips25_sap3/_0659_ sg13g2_a221oi_1
XFILLER_32_146 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3077_ heichips25_sap3/_0690_ heichips25_sap3/net249 heichips25_sap3/_1668_
+ VPWR VGND sg13g2_nand2b_1
Xheichips25_sap3__2028_ heichips25_sap3/net259 heichips25_sap3/_1361_ heichips25_sap3/_1449_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_can_lehmann_fsm_fanout407 heichips25_can_lehmann_fsm/net408 heichips25_can_lehmann_fsm/net407
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout429 heichips25_can_lehmann_fsm/net431 heichips25_can_lehmann_fsm/net429
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout418 heichips25_can_lehmann_fsm/net419 heichips25_can_lehmann_fsm/net418
+ VPWR VGND sg13g2_buf_1
Xheichips25_sap3__3979_ heichips25_sap3/net443 VGND VPWR heichips25_sap3/_0120_ heichips25_sap3__3979_/Q
+ clkload19/A sg13g2_dfrbpq_1
XFILLER_28_408 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2703_ VGND VPWR heichips25_can_lehmann_fsm/_0869_ heichips25_can_lehmann_fsm/net385
+ heichips25_can_lehmann_fsm/_0251_ heichips25_can_lehmann_fsm/_0817_ sg13g2_a21oi_1
Xclkbuf_5_12__f_heichips25_sap3\_sap_3_inst.alu_inst.clk heichips25_sap3__4009_/CLK
+ clknet_4_6_0_heichips25_sap3\/sap_3_inst.alu_inst.clk VPWR VGND sg13g2_buf_16
XFILLER_23_113 VPWR VGND sg13g2_fill_2
XFILLER_24_614 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2634_ heichips25_can_lehmann_fsm/net465 VPWR heichips25_can_lehmann_fsm/_0783_
+ VGND heichips25_can_lehmann_fsm/net964 heichips25_can_lehmann_fsm/net394 sg13g2_o21ai_1
XFILLER_23_124 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2565_ VGND VPWR heichips25_can_lehmann_fsm/_0906_ heichips25_can_lehmann_fsm/net377
+ heichips25_can_lehmann_fsm/_0182_ heichips25_can_lehmann_fsm/_0748_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2496_ heichips25_can_lehmann_fsm/net467 VPWR heichips25_can_lehmann_fsm/_0714_
+ VGND heichips25_can_lehmann_fsm/net962 heichips25_can_lehmann_fsm/net355 sg13g2_o21ai_1
XFILLER_3_518 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__3048_ net605 VGND VPWR heichips25_can_lehmann_fsm/_0273_
+ heichips25_can_lehmann_fsm__3048_/Q clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_36_76 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3000_ heichips25_sap3/_0627_ net44 heichips25_sap3/net201 VPWR VGND
+ sg13g2_nand2_1
XFILLER_15_625 VPWR VGND sg13g2_fill_2
XFILLER_14_135 VPWR VGND sg13g2_decap_4
XFILLER_15_669 VPWR VGND sg13g2_decap_4
XFILLER_14_179 VPWR VGND sg13g2_fill_2
XFILLER_23_680 VPWR VGND sg13g2_fill_1
Xinput18 uio_in[7] net18 VPWR VGND sg13g2_buf_1
XFILLER_7_802 VPWR VGND sg13g2_fill_1
XFILLER_22_190 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3902_ heichips25_sap3/net449 VGND VPWR heichips25_sap3/_0043_ heichips25_sap3__3902_/Q
+ heichips25_sap3__3920_/CLK sg13g2_dfrbpq_1
Xheichips25_sap3__3833_ VGND VPWR heichips25_sap3__3970_/Q heichips25_sap3/_1279_
+ heichips25_sap3/_1338_ heichips25_sap3/net291 sg13g2_a21oi_1
Xheichips25_sap3__3764_ heichips25_sap3__4042_/Q heichips25_sap3__4043_/Q heichips25_sap3/_1275_
+ heichips25_sap3/_1276_ VPWR VGND sg13g2_a21o_1
Xheichips25_sap3__3695_ heichips25_sap3/_0150_ heichips25_sap3/_1194_ heichips25_sap3/_1229_
+ heichips25_sap3/net113 heichips25_sap3/_1414_ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2715_ heichips25_sap3__3917_/Q heichips25_sap3/net284 heichips25_sap3/_0361_
+ VPWR VGND sg13g2_xor2_1
Xheichips25_sap3__2646_ heichips25_sap3/_1719_ heichips25_sap3/_0312_ heichips25_sap3/_0313_
+ VPWR VGND sg13g2_and2_1
XFILLER_38_717 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2577_ heichips25_sap3/_1680_ heichips25_sap3/_1713_ heichips25_sap3__3973_/Q
+ heichips25_sap3/_0250_ VPWR VGND heichips25_sap3/_1731_ sg13g2_nand4_1
XFILLER_18_452 VPWR VGND sg13g2_fill_1
XFILLER_46_783 VPWR VGND sg13g2_fill_2
XFILLER_45_271 VPWR VGND sg13g2_fill_1
XFILLER_19_997 VPWR VGND sg13g2_fill_2
XFILLER_33_400 VPWR VGND sg13g2_decap_4
XFILLER_34_989 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3129_ heichips25_sap3/_0738_ heichips25_sap3/_0739_ heichips25_sap3/_0741_
+ heichips25_sap3/_0742_ VPWR VGND sg13g2_nor3_1
Xheichips25_can_lehmann_fsm__2350_ heichips25_can_lehmann_fsm/net494 VPWR heichips25_can_lehmann_fsm/_0641_
+ VGND heichips25_can_lehmann_fsm/net857 heichips25_can_lehmann_fsm/net423 sg13g2_o21ai_1
XFILLER_14_680 VPWR VGND sg13g2_decap_8
XFILLER_9_161 VPWR VGND sg13g2_fill_2
XFILLER_20_149 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2281_ heichips25_can_lehmann_fsm/net1170 VPWR heichips25_can_lehmann_fsm/_0595_
+ VGND heichips25_can_lehmann_fsm__2826_/Q heichips25_can_lehmann_fsm/_1047_ sg13g2_o21ai_1
XFILLER_29_717 VPWR VGND sg13g2_fill_1
XFILLER_28_227 VPWR VGND sg13g2_fill_2
XFILLER_44_709 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__1996_ heichips25_can_lehmann_fsm/_0352_ heichips25_can_lehmann_fsm/net185
+ heichips25_can_lehmann_fsm/_0351_ VPWR VGND sg13g2_nand2_1
XFILLER_43_219 VPWR VGND sg13g2_fill_1
XFILLER_25_934 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2617_ VGND VPWR heichips25_can_lehmann_fsm/_0893_ heichips25_can_lehmann_fsm/net373
+ heichips25_can_lehmann_fsm/_0208_ heichips25_can_lehmann_fsm/_0774_ sg13g2_a21oi_1
XFILLER_24_455 VPWR VGND sg13g2_fill_1
XFILLER_7_109 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2548_ heichips25_can_lehmann_fsm/net473 VPWR heichips25_can_lehmann_fsm/_0740_
+ VGND heichips25_can_lehmann_fsm/net1037 heichips25_can_lehmann_fsm/net364 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2479_ VGND VPWR heichips25_can_lehmann_fsm/_0928_ heichips25_can_lehmann_fsm/net416
+ heichips25_can_lehmann_fsm/_0139_ heichips25_can_lehmann_fsm/_0705_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__3031__614 VPWR VGND net613 sg13g2_tiehi
Xheichips25_sap3__3480_ heichips25_sap3/_0863_ heichips25_sap3/_1021_ heichips25_sap3/_1079_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__2500_ heichips25_sap3/_1913_ heichips25_sap3/_1909_ heichips25_sap3/_1912_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__2431_ heichips25_sap3/_1846_ heichips25_sap3/net75 heichips25_sap3__3983_/Q
+ heichips25_sap3/net81 heichips25_sap3__3967_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2362_ heichips25_sap3/_1783_ heichips25_sap3/_1472_ heichips25_sap3/_1496_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__2293_ heichips25_sap3/net227 heichips25_sap3/_1613_ heichips25_sap3/net273
+ heichips25_sap3/_1714_ VPWR VGND sg13g2_nand3_1
XFILLER_28_783 VPWR VGND sg13g2_fill_2
XFILLER_34_208 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__4032_ heichips25_sap3/net458 VGND VPWR heichips25_sap3/_0173_ heichips25_sap3__4032_/Q
+ clknet_leaf_1_clk sg13g2_dfrbpq_1
XFILLER_30_403 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2825__557 VPWR VGND net556 sg13g2_tiehi
XFILLER_42_296 VPWR VGND sg13g2_decap_8
XFILLER_8_25 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm_hold871 heichips25_can_lehmann_fsm__2889_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net870 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold860 heichips25_can_lehmann_fsm/_0154_ VPWR VGND heichips25_can_lehmann_fsm/net859
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold882 heichips25_can_lehmann_fsm__3011_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net881 sg13g2_dlygate4sd3_1
XFILLER_6_175 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3816_ heichips25_sap3/_1323_ heichips25_sap3/_1278_ heichips25_sap3__4008_/Q
+ heichips25_sap3/_1272_ heichips25_sap3__3976_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3747_ heichips25_sap3/_1257_ heichips25_sap3/_1258_ heichips25_sap3/_1259_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__3678_ heichips25_sap3/_1036_ heichips25_sap3/_1017_ heichips25_sap3/_1220_
+ VPWR VGND sg13g2_xor2_1
Xheichips25_sap3__2629_ heichips25_sap3/_1559_ VPWR heichips25_sap3/_0296_ VGND heichips25_sap3/_1522_
+ heichips25_sap3/_1526_ sg13g2_o21ai_1
X_15_ net516 uio_out_sap3\[1\] net504 net28 VPWR VGND sg13g2_mux2_1
XFILLER_19_750 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1850_ heichips25_can_lehmann_fsm/_1139_ heichips25_can_lehmann_fsm/_1162_
+ heichips25_can_lehmann_fsm/_1166_ VPWR VGND sg13g2_nor2_1
Xheichips25_can_lehmann_fsm__1781_ heichips25_can_lehmann_fsm/net1215 heichips25_can_lehmann_fsm__2803_/Q
+ heichips25_can_lehmann_fsm__2802_/Q heichips25_can_lehmann_fsm/_1097_ VPWR VGND
+ sg13g2_nor3_1
Xheichips25_sap3_fanout119 heichips25_sap3/_0750_ heichips25_sap3/net119 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout108 heichips25_sap3/net110 heichips25_sap3/net108 VPWR VGND
+ sg13g2_buf_1
Xheichips25_can_lehmann_fsm_hold1209 heichips25_can_lehmann_fsm/_0037_ VPWR VGND heichips25_can_lehmann_fsm/net1208
+ sg13g2_dlygate4sd3_1
XFILLER_21_414 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2402_ heichips25_can_lehmann_fsm/net473 VPWR heichips25_can_lehmann_fsm/_0667_
+ VGND heichips25_can_lehmann_fsm__2875_/Q heichips25_can_lehmann_fsm/net364 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2333_ VGND VPWR heichips25_can_lehmann_fsm/_0968_ heichips25_can_lehmann_fsm/net363
+ heichips25_can_lehmann_fsm/_0066_ heichips25_can_lehmann_fsm/_0632_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2264_ heichips25_can_lehmann_fsm/net327 VPWR heichips25_can_lehmann_fsm/_0582_
+ VGND heichips25_can_lehmann_fsm/net1181 heichips25_can_lehmann_fsm/net208 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__3058__783 VPWR VGND net782 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2195_ VGND VPWR heichips25_can_lehmann_fsm/_0525_ heichips25_can_lehmann_fsm/_0526_
+ heichips25_can_lehmann_fsm/_0033_ heichips25_can_lehmann_fsm/_0527_ sg13g2_a21oi_1
XFILLER_29_514 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1979_ heichips25_can_lehmann_fsm/net323 VPWR heichips25_can_lehmann_fsm/_0338_
+ VGND heichips25_can_lehmann_fsm/net1257 heichips25_can_lehmann_fsm/net179 sg13g2_o21ai_1
XFILLER_40_701 VPWR VGND sg13g2_fill_1
XFILLER_25_764 VPWR VGND sg13g2_decap_4
XFILLER_25_775 VPWR VGND sg13g2_fill_1
XFILLER_33_11 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2980_ heichips25_sap3/_0614_ heichips25_sap3__3910_/Q heichips25_sap3/_0607_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__3601_ VPWR heichips25_sap3/_0112_ heichips25_sap3/_1173_ VGND sg13g2_inv_1
Xheichips25_sap3__3532_ heichips25_sap3/net120 heichips25_sap3/_1024_ heichips25_sap3/_1123_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_can_lehmann_fsm__2935__596 VPWR VGND net595 sg13g2_tiehi
Xheichips25_sap3__3463_ heichips25_sap3/_1064_ heichips25_sap3/_1065_ heichips25_sap3/_0933_
+ heichips25_sap3/_1066_ VPWR VGND sg13g2_nand3_1
Xheichips25_sap3__2414_ VPWR VGND heichips25_sap3/_1830_ heichips25_sap3/_1654_ heichips25_sap3/_1827_
+ heichips25_sap3/_1404_ heichips25_sap3/_1831_ heichips25_sap3/net91 sg13g2_a221oi_1
Xheichips25_sap3__3394_ heichips25_sap3/_0802_ VPWR heichips25_sap3/_1002_ VGND heichips25_sap3/net63
+ heichips25_sap3/_0855_ sg13g2_o21ai_1
XFILLER_47_388 VPWR VGND sg13g2_fill_2
XFILLER_35_528 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2345_ heichips25_sap3/_1765_ VPWR heichips25_sap3/_1766_ VGND heichips25_sap3/_1756_
+ heichips25_sap3/_1764_ sg13g2_o21ai_1
Xheichips25_sap3__2276_ VGND VPWR heichips25_sap3/net234 heichips25_sap3/net225 heichips25_sap3/_1697_
+ heichips25_sap3/_1516_ sg13g2_a21oi_1
XFILLER_15_241 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__4015_ heichips25_sap3/net439 VGND VPWR heichips25_sap3/_0156_ heichips25_sap3__4015_/Q
+ heichips25_sap3__4015_/CLK sg13g2_dfrbpq_1
XFILLER_15_274 VPWR VGND sg13g2_fill_1
XFILLER_31_734 VPWR VGND sg13g2_fill_1
XFILLER_8_952 VPWR VGND sg13g2_decap_8
XFILLER_8_963 VPWR VGND sg13g2_fill_1
XFILLER_7_462 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2877__742 VPWR VGND net741 sg13g2_tiehi
XFILLER_7_495 VPWR VGND sg13g2_decap_4
XFILLER_48_1021 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2951_ net531 VGND VPWR heichips25_can_lehmann_fsm/net1078
+ heichips25_can_lehmann_fsm__2951_/Q clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_38_322 VPWR VGND sg13g2_decap_8
XFILLER_38_300 VPWR VGND sg13g2_fill_2
XFILLER_39_878 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2882_ net731 VGND VPWR heichips25_can_lehmann_fsm/_0107_
+ heichips25_can_lehmann_fsm__2882_/Q clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_17_0 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1902_ VGND VPWR heichips25_can_lehmann_fsm/_1205_ heichips25_can_lehmann_fsm/_1206_
+ heichips25_can_lehmann_fsm/_1215_ heichips25_can_lehmann_fsm/_1214_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__1833_ heichips25_can_lehmann_fsm/_1148_ VPWR heichips25_can_lehmann_fsm/_1149_
+ VGND heichips25_can_lehmann_fsm/net343 heichips25_can_lehmann_fsm/_0985_ sg13g2_o21ai_1
XFILLER_41_509 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1764_ uo_out_fsm\[6\] heichips25_can_lehmann_fsm/_1080_
+ heichips25_can_lehmann_fsm/_1081_ VPWR VGND sg13g2_nand2_1
Xheichips25_can_lehmann_fsm_hold1028 heichips25_can_lehmann_fsm__2955_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1027 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1006 heichips25_can_lehmann_fsm__2940_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1005 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__1695_ heichips25_can_lehmann_fsm/_1019_ heichips25_can_lehmann_fsm/net305
+ heichips25_can_lehmann_fsm__2944_/Q heichips25_can_lehmann_fsm/net313 heichips25_can_lehmann_fsm__2920_/Q
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm_hold1039 heichips25_can_lehmann_fsm__2962_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1038 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1017 heichips25_can_lehmann_fsm/_0100_ VPWR VGND heichips25_can_lehmann_fsm/net1016
+ sg13g2_dlygate4sd3_1
XFILLER_21_222 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2316_ net8 net9 heichips25_can_lehmann_fsm/_0623_ VPWR
+ VGND sg13g2_and2_1
Xheichips25_can_lehmann_fsm__2247_ VGND VPWR heichips25_can_lehmann_fsm/net911 heichips25_can_lehmann_fsm/net170
+ heichips25_can_lehmann_fsm/_0568_ heichips25_can_lehmann_fsm/_0567_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2778__651 VPWR VGND net650 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2178_ heichips25_can_lehmann_fsm/net325 VPWR heichips25_can_lehmann_fsm/_0514_
+ VGND heichips25_can_lehmann_fsm/net1202 heichips25_can_lehmann_fsm/net160 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2971__741 VPWR VGND net740 sg13g2_tiehi
XFILLER_0_159 VPWR VGND sg13g2_fill_2
XFILLER_28_44 VPWR VGND sg13g2_decap_4
XFILLER_28_55 VPWR VGND sg13g2_fill_1
XFILLER_44_314 VPWR VGND sg13g2_fill_1
XFILLER_44_32 VPWR VGND sg13g2_decap_8
Xheichips25_sap3_fanout450 heichips25_sap3/net463 heichips25_sap3/net450 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3__2130_ heichips25_sap3/net251 heichips25_sap3/net250 heichips25_sap3/_1551_
+ VPWR VGND sg13g2_and2_1
Xheichips25_sap3_fanout461 heichips25_sap3/net462 heichips25_sap3/net461 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3__2061_ heichips25_sap3/_1476_ heichips25_sap3/_1481_ heichips25_sap3/_1482_
+ VPWR VGND sg13g2_and2_1
Xheichips25_sap3_hold1072 heichips25_sap3__4046_/Q VPWR VGND heichips25_sap3/net1071
+ sg13g2_dlygate4sd3_1
XFILLER_12_244 VPWR VGND sg13g2_decap_8
XFILLER_8_237 VPWR VGND sg13g2_fill_2
XFILLER_8_259 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2963_ VGND VPWR heichips25_sap3/net65 heichips25_sap3/_0588_ heichips25_sap3/_0601_
+ heichips25_sap3/_0436_ sg13g2_a21oi_1
XFILLER_5_37 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2894_ VGND VPWR heichips25_sap3/net65 heichips25_sap3/_0522_ heichips25_sap3/_0535_
+ heichips25_sap3/net203 sg13g2_a21oi_1
Xheichips25_sap3__3515_ heichips25_sap3/net106 heichips25_sap3/_1108_ heichips25_sap3/_1109_
+ VPWR VGND sg13g2_nor2_1
XFILLER_48_653 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3446_ heichips25_sap3/_0079_ heichips25_sap3/_1041_ heichips25_sap3/_1051_
+ heichips25_sap3/_0748_ heichips25_sap3/_1420_ VPWR VGND sg13g2_a22oi_1
XFILLER_35_314 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3377_ VPWR VGND heichips25_sap3__4000_/Q heichips25_sap3/net124
+ heichips25_sap3/net146 heichips25_sap3__4016_/Q heichips25_sap3/_0985_ heichips25_sap3/net116
+ sg13g2_a221oi_1
Xheichips25_sap3__2328_ heichips25_sap3/_1749_ heichips25_sap3/net79 heichips25_sap3__4026_/Q
+ heichips25_sap3/net81 heichips25_sap3__3970_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2259_ heichips25_sap3/_1456_ heichips25_sap3/_1677_ heichips25_sap3/_1678_
+ heichips25_sap3/_1679_ heichips25_sap3/_1680_ VPWR VGND sg13g2_and4_1
Xheichips25_can_lehmann_fsm__2101_ heichips25_can_lehmann_fsm/_0441_ heichips25_can_lehmann_fsm/net344
+ heichips25_can_lehmann_fsm/net200 VPWR VGND sg13g2_nand2_1
Xclkbuf_4_11_0_heichips25_sap3\_sap_3_inst.alu_inst.clk clknet_0_heichips25_sap3\/sap_3_inst.alu_inst.clk
+ clknet_4_11_0_heichips25_sap3\/sap_3_inst.alu_inst.clk VPWR VGND sg13g2_buf_8
Xheichips25_can_lehmann_fsm__2032_ heichips25_can_lehmann_fsm/net324 VPWR heichips25_can_lehmann_fsm/_0383_
+ VGND heichips25_can_lehmann_fsm/net1244 heichips25_can_lehmann_fsm/net177 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2934_ net599 VGND VPWR heichips25_can_lehmann_fsm/net864
+ heichips25_can_lehmann_fsm__2934_/Q clknet_leaf_14_clk sg13g2_dfrbpq_1
XFILLER_39_664 VPWR VGND sg13g2_fill_2
XFILLER_38_163 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2865_ net765 VGND VPWR heichips25_can_lehmann_fsm/net884
+ heichips25_can_lehmann_fsm__2865_/Q clknet_leaf_8_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2796_ net614 VGND VPWR heichips25_can_lehmann_fsm/_0021_
+ heichips25_can_lehmann_fsm__2796_/Q clknet_leaf_3_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1816_ heichips25_can_lehmann_fsm/_0985_ heichips25_can_lehmann_fsm/_0987_
+ heichips25_can_lehmann_fsm/_1122_ heichips25_can_lehmann_fsm/_1132_ VPWR VGND sg13g2_mux2_1
Xheichips25_can_lehmann_fsm__1747_ heichips25_can_lehmann_fsm/_1064_ heichips25_can_lehmann_fsm/_1066_
+ heichips25_can_lehmann_fsm/_1061_ heichips25_can_lehmann_fsm/_1067_ VPWR VGND sg13g2_nand3_1
XFILLER_14_24 VPWR VGND sg13g2_decap_8
XFILLER_22_553 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1678_ heichips25_can_lehmann_fsm/net338 heichips25_can_lehmann_fsm/_0989_
+ heichips25_can_lehmann_fsm/_1002_ VPWR VGND sg13g2_and2_1
Xheichips25_sap3__3881__826 VPWR net825 heichips25_sap3__4013_/CLK VGND sg13g2_inv_1
XFILLER_2_903 VPWR VGND sg13g2_fill_1
XFILLER_2_958 VPWR VGND sg13g2_decap_8
XFILLER_39_98 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3300_ VGND VPWR heichips25_sap3/net127 heichips25_sap3/_0911_ heichips25_sap3/_0912_
+ heichips25_sap3/_0863_ sg13g2_a21oi_1
Xheichips25_sap3__3231_ heichips25_sap3/_0844_ heichips25_sap3__3972_/Q heichips25_sap3/net134
+ VPWR VGND sg13g2_nand2_1
XFILLER_45_656 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3162_ heichips25_sap3/_0761_ heichips25_sap3/_0765_ heichips25_sap3/_0756_
+ heichips25_sap3/_0775_ VPWR VGND heichips25_sap3/_0774_ sg13g2_nand4_1
Xheichips25_sap3__2113_ heichips25_sap3/_1528_ heichips25_sap3/_1533_ heichips25_sap3/_1534_
+ VPWR VGND sg13g2_and2_1
XFILLER_26_892 VPWR VGND sg13g2_fill_1
XFILLER_32_306 VPWR VGND sg13g2_decap_8
Xheichips25_sap3_fanout291 heichips25_sap3/_1276_ heichips25_sap3/net291 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3__3093_ heichips25_sap3/_1530_ heichips25_sap3/_1544_ heichips25_sap3/net271
+ heichips25_sap3/_0706_ VPWR VGND heichips25_sap3/_0705_ sg13g2_nand4_1
Xheichips25_sap3_fanout280 heichips25_sap3__3903_/Q heichips25_sap3/net280 VPWR VGND
+ sg13g2_buf_1
XFILLER_41_895 VPWR VGND sg13g2_fill_2
XFILLER_40_372 VPWR VGND sg13g2_fill_1
XFILLER_40_350 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2044_ heichips25_sap3__4064_/Q heichips25_sap3/_1458_ heichips25_sap3/_1465_
+ VPWR VGND sg13g2_nor2_1
XFILLER_5_730 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3995_ heichips25_sap3/net439 VGND VPWR heichips25_sap3/_0136_ heichips25_sap3__3995_/Q
+ heichips25_sap3__4015_/CLK sg13g2_dfrbpq_1
Xheichips25_sap3__2946_ net47 heichips25_sap3/_0434_ heichips25_sap3/_0584_ VPWR VGND
+ sg13g2_nor2b_1
XFILLER_45_1002 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2877_ net46 heichips25_sap3/net157 heichips25_sap3/_0518_ VPWR VGND
+ sg13g2_nor2b_1
Xheichips25_sap3__3429_ heichips25_sap3/_1031_ heichips25_sap3/_1032_ heichips25_sap3/_1033_
+ heichips25_sap3/_1034_ heichips25_sap3/_1035_ VPWR VGND sg13g2_and4_1
XFILLER_36_678 VPWR VGND sg13g2_decap_4
XFILLER_24_807 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2650_ heichips25_can_lehmann_fsm/net491 VPWR heichips25_can_lehmann_fsm/_0791_
+ VGND heichips25_can_lehmann_fsm__3000_/Q heichips25_can_lehmann_fsm/net421 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__1601_ VPWR heichips25_can_lehmann_fsm/_0925_ heichips25_can_lehmann_fsm/net981
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__2581_ VGND VPWR heichips25_can_lehmann_fsm/_0902_ heichips25_can_lehmann_fsm/net369
+ heichips25_can_lehmann_fsm/_0190_ heichips25_can_lehmann_fsm/_0756_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__1532_ VPWR heichips25_can_lehmann_fsm/_0856_ heichips25_can_lehmann_fsm/net1155
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__2015_ VGND VPWR heichips25_can_lehmann_fsm/net178 heichips25_can_lehmann_fsm/_0367_
+ heichips25_can_lehmann_fsm/_0012_ heichips25_can_lehmann_fsm/_0368_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2917_ net661 VGND VPWR heichips25_can_lehmann_fsm/_0142_
+ heichips25_can_lehmann_fsm__2917_/Q clknet_leaf_18_clk sg13g2_dfrbpq_1
XFILLER_26_111 VPWR VGND sg13g2_fill_2
XFILLER_27_623 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2848_ net799 VGND VPWR heichips25_can_lehmann_fsm/_0073_
+ heichips25_can_lehmann_fsm__2848_/Q clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_41_136 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2779_ net648 VGND VPWR heichips25_can_lehmann_fsm/net1254
+ heichips25_can_lehmann_fsm__2779_/Q clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_10_501 VPWR VGND sg13g2_decap_4
XFILLER_22_372 VPWR VGND sg13g2_fill_2
XFILLER_23_895 VPWR VGND sg13g2_fill_2
XFILLER_10_545 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2903__690 VPWR VGND net689 sg13g2_tiehi
Xheichips25_sap3__2800_ heichips25_sap3/_1885_ heichips25_sap3/net169 heichips25_sap3/_0445_
+ VPWR VGND sg13g2_nor2b_1
Xheichips25_sap3__3780_ heichips25_sap3/_1291_ heichips25_sap3/_1274_ heichips25_sap3__3940_/Q
+ heichips25_sap3/_1270_ heichips25_sap3__4020_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2731_ heichips25_sap3/_0357_ heichips25_sap3/_0359_ heichips25_sap3/_0377_
+ VPWR VGND sg13g2_and2_1
XFILLER_2_755 VPWR VGND sg13g2_fill_1
XFILLER_2_744 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2662_ heichips25_sap3/_0326_ heichips25_sap3__4066_/Q heichips25_sap3/_1554_
+ VPWR VGND sg13g2_nand2_1
XFILLER_1_276 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2593_ heichips25_sap3/_0266_ heichips25_sap3/net86 heichips25_sap3__3957_/Q
+ heichips25_sap3/net89 heichips25_sap3__3941_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3214_ heichips25_sap3/_0827_ heichips25_sap3__3955_/Q heichips25_sap3/net108
+ VPWR VGND sg13g2_nand2_1
XFILLER_17_177 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3145_ heichips25_sap3/_0758_ heichips25_sap3/net152 heichips25_sap3/net150
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__3076_ heichips25_sap3/_1462_ heichips25_sap3/_1508_ heichips25_sap3/_0689_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__2027_ heichips25_sap3/net269 heichips25_sap3/net268 heichips25_sap3/_1448_
+ VPWR VGND heichips25_sap3/net273 sg13g2_nand3b_1
XFILLER_9_365 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3978_ heichips25_sap3/net444 VGND VPWR heichips25_sap3/_0119_ heichips25_sap3__3978_/Q
+ clkload21/A sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm_fanout408 heichips25_can_lehmann_fsm/net432 heichips25_can_lehmann_fsm/net408
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout419 heichips25_can_lehmann_fsm/net420 heichips25_can_lehmann_fsm/net419
+ VPWR VGND sg13g2_buf_1
Xheichips25_sap3__2929_ heichips25_sap3/_0568_ heichips25_sap3/_0350_ heichips25_sap3/_0445_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_can_lehmann_fsm__2835__537 VPWR VGND net536 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__3052__767 VPWR VGND net766 sg13g2_tiehi
XFILLER_48_291 VPWR VGND sg13g2_fill_2
XFILLER_37_954 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2702_ heichips25_can_lehmann_fsm/net497 VPWR heichips25_can_lehmann_fsm/_0817_
+ VGND heichips25_can_lehmann_fsm/net1076 heichips25_can_lehmann_fsm/net385 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2633_ VGND VPWR heichips25_can_lehmann_fsm/_0889_ heichips25_can_lehmann_fsm/net361
+ heichips25_can_lehmann_fsm/_0216_ heichips25_can_lehmann_fsm/_0782_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2564_ heichips25_can_lehmann_fsm/net488 VPWR heichips25_can_lehmann_fsm/_0748_
+ VGND heichips25_can_lehmann_fsm__2956_/Q heichips25_can_lehmann_fsm/net377 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2495_ VGND VPWR heichips25_can_lehmann_fsm/_0924_ heichips25_can_lehmann_fsm/net390
+ heichips25_can_lehmann_fsm/_0147_ heichips25_can_lehmann_fsm/_0713_ sg13g2_a21oi_1
XFILLER_31_191 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__3047_ net637 VGND VPWR heichips25_can_lehmann_fsm/_0272_
+ heichips25_can_lehmann_fsm__3047_/Q clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_36_55 VPWR VGND sg13g2_fill_1
XFILLER_27_431 VPWR VGND sg13g2_decap_8
XFILLER_36_99 VPWR VGND sg13g2_fill_2
XFILLER_14_158 VPWR VGND sg13g2_decap_8
XFILLER_7_825 VPWR VGND sg13g2_fill_1
XFILLER_6_302 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3901_ heichips25_sap3/net448 VGND VPWR heichips25_sap3/_0042_ heichips25_sap3__3901_/Q
+ clkload24/A sg13g2_dfrbpq_1
XFILLER_6_324 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3832_ heichips25_sap3/_1337_ heichips25_sap3/_1265_ heichips25_sap3__4002_/Q
+ heichips25_sap3/_1259_ heichips25_sap3__3986_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_6_368 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3763_ heichips25_sap3__4040_/Q heichips25_sap3__4041_/Q heichips25_sap3__4043_/Q
+ heichips25_sap3__4042_/Q heichips25_sap3/_1275_ VPWR VGND sg13g2_nor4_1
Xheichips25_sap3__2714_ heichips25_sap3/net284 heichips25_sap3__3917_/Q heichips25_sap3/_0360_
+ VPWR VGND sg13g2_and2_1
Xheichips25_sap3__3694_ heichips25_sap3/net111 heichips25_sap3/_1079_ heichips25_sap3/_1229_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__2645_ heichips25_sap3/_0312_ heichips25_sap3/_1623_ heichips25_sap3/net230
+ heichips25_sap3/_1605_ heichips25_sap3/_1476_ VPWR VGND sg13g2_a22oi_1
XFILLER_38_707 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2576_ heichips25_sap3/_1695_ heichips25_sap3/_1713_ heichips25_sap3__3941_/Q
+ heichips25_sap3/_0249_ VPWR VGND heichips25_sap3/_1731_ sg13g2_nand4_1
XFILLER_18_431 VPWR VGND sg13g2_fill_1
XFILLER_19_965 VPWR VGND sg13g2_fill_1
XFILLER_19_976 VPWR VGND sg13g2_fill_1
XFILLER_45_250 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3128_ heichips25_sap3/_1758_ heichips25_sap3/_0740_ heichips25_sap3/_1659_
+ heichips25_sap3/_0741_ VPWR VGND sg13g2_nand3_1
XFILLER_13_191 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3059_ heichips25_sap3/net239 heichips25_sap3/_1721_ heichips25_sap3/_1449_
+ heichips25_sap3/_0672_ VPWR VGND sg13g2_nand3_1
Xheichips25_can_lehmann_fsm__2280_ VGND VPWR heichips25_can_lehmann_fsm/net208 heichips25_can_lehmann_fsm/_0593_
+ heichips25_can_lehmann_fsm/_0051_ heichips25_can_lehmann_fsm/_0594_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm_fanout205 heichips25_can_lehmann_fsm/net210 heichips25_can_lehmann_fsm/net205
+ VPWR VGND sg13g2_buf_1
XFILLER_47_0 VPWR VGND sg13g2_fill_2
XFILLER_3_81 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2887__722 VPWR VGND net721 sg13g2_tiehi
XFILLER_28_206 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1995_ heichips25_can_lehmann_fsm/_0351_ heichips25_can_lehmann_fsm__2785_/Q
+ heichips25_can_lehmann_fsm/_1067_ VPWR VGND sg13g2_xnor2_1
XFILLER_43_209 VPWR VGND sg13g2_fill_1
XFILLER_36_272 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2616_ heichips25_can_lehmann_fsm/net486 VPWR heichips25_can_lehmann_fsm/_0774_
+ VGND heichips25_can_lehmann_fsm__2982_/Q heichips25_can_lehmann_fsm/net373 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2547_ VGND VPWR heichips25_can_lehmann_fsm/_0911_ heichips25_can_lehmann_fsm/net392
+ heichips25_can_lehmann_fsm/_0173_ heichips25_can_lehmann_fsm/_0739_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2478_ heichips25_can_lehmann_fsm/net483 VPWR heichips25_can_lehmann_fsm/_0705_
+ VGND heichips25_can_lehmann_fsm/net869 heichips25_can_lehmann_fsm/net416 sg13g2_o21ai_1
XFILLER_22_35 VPWR VGND sg13g2_decap_8
XFILLER_3_327 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2430_ heichips25_sap3/_1845_ heichips25_sap3/net85 heichips25_sap3__3951_/Q
+ heichips25_sap3/net87 heichips25_sap3__3943_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2361_ heichips25_sap3/_1458_ heichips25_sap3/_1460_ heichips25_sap3/_1613_
+ heichips25_sap3/_1782_ VPWR VGND sg13g2_nor3_1
Xheichips25_can_lehmann_fsm__2788__631 VPWR VGND net630 sg13g2_tiehi
Xheichips25_sap3__2292_ heichips25_sap3/_1708_ heichips25_sap3/_1707_ heichips25_sap3/_1711_
+ heichips25_sap3/_1713_ VPWR VGND sg13g2_a21o_1
Xheichips25_sap3__4031_ heichips25_sap3/net461 VGND VPWR heichips25_sap3/net837 heichips25_sap3__4031_/Q
+ clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_42_264 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm_hold850 heichips25_can_lehmann_fsm__3022_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net849 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold861 heichips25_can_lehmann_fsm__2998_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net860 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold883 heichips25_can_lehmann_fsm/_0236_ VPWR VGND heichips25_can_lehmann_fsm/net882
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold872 heichips25_can_lehmann_fsm/_0114_ VPWR VGND heichips25_can_lehmann_fsm/net871
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold894 heichips25_can_lehmann_fsm__2923_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net893 sg13g2_dlygate4sd3_1
XFILLER_6_132 VPWR VGND sg13g2_decap_8
XFILLER_10_183 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3815_ heichips25_sap3/_1322_ heichips25_sap3/_1281_ heichips25_sap3__4016_/Q
+ heichips25_sap3/_1279_ heichips25_sap3__3968_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3746_ heichips25_sap3/_1258_ heichips25_sap3/_1428_ heichips25_sap3__4041_/Q
+ VPWR VGND sg13g2_nand2_1
XFILLER_3_883 VPWR VGND sg13g2_fill_2
XFILLER_3_850 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3677_ heichips25_sap3/_0142_ heichips25_sap3/_1122_ heichips25_sap3/_1219_
+ heichips25_sap3/net111 heichips25_sap3/_1415_ VPWR VGND sg13g2_a22oi_1
XFILLER_2_382 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2628_ heichips25_sap3/_1435_ heichips25_sap3/_1448_ heichips25_sap3/_1464_
+ heichips25_sap3/_1478_ heichips25_sap3/_0295_ VPWR VGND sg13g2_nor4_1
X_14_ net515 uio_out_sap3\[0\] net504 net27 VPWR VGND sg13g2_mux2_1
Xheichips25_sap3__2559_ heichips25_sap3/_0233_ VPWR heichips25_sap3/_0234_ VGND heichips25_sap3/_1367_
+ heichips25_sap3/net155 sg13g2_o21ai_1
Xheichips25_sap3_fanout109 heichips25_sap3/net110 heichips25_sap3/net109 VPWR VGND
+ sg13g2_buf_1
Xheichips25_can_lehmann_fsm__1780_ heichips25_can_lehmann_fsm/_1095_ VPWR heichips25_can_lehmann_fsm/_1096_
+ VGND heichips25_can_lehmann_fsm__2869_/Q heichips25_can_lehmann_fsm/net335 sg13g2_o21ai_1
XFILLER_34_765 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2401_ VGND VPWR heichips25_can_lehmann_fsm/_0951_ heichips25_can_lehmann_fsm/net390
+ heichips25_can_lehmann_fsm/_0100_ heichips25_can_lehmann_fsm/_0666_ sg13g2_a21oi_1
XFILLER_33_275 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2332_ heichips25_can_lehmann_fsm/net475 VPWR heichips25_can_lehmann_fsm/_0632_
+ VGND heichips25_can_lehmann_fsm__2840_/Q heichips25_can_lehmann_fsm/net363 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2263_ VGND VPWR heichips25_can_lehmann_fsm/net939 heichips25_can_lehmann_fsm/net173
+ heichips25_can_lehmann_fsm/_0581_ heichips25_can_lehmann_fsm/_0580_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2194_ heichips25_can_lehmann_fsm/net325 VPWR heichips25_can_lehmann_fsm/_0527_
+ VGND heichips25_can_lehmann_fsm/net1192 heichips25_can_lehmann_fsm/net160 sg13g2_o21ai_1
Xclkbuf_5_13__f_heichips25_sap3\_sap_3_inst.alu_inst.clk clkload21/A clknet_4_6_0_heichips25_sap3\/sap_3_inst.alu_inst.clk
+ VPWR VGND sg13g2_buf_16
XFILLER_44_518 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__1978_ heichips25_can_lehmann_fsm__2799_/Q heichips25_can_lehmann_fsm/net183
+ heichips25_can_lehmann_fsm/_0337_ VPWR VGND sg13g2_nor2_1
XFILLER_24_275 VPWR VGND sg13g2_decap_8
XFILLER_25_787 VPWR VGND sg13g2_fill_2
XFILLER_33_23 VPWR VGND sg13g2_fill_1
Xheichips25_sap3_hold1276 heichips25_sap3__4029_/Q VPWR VGND heichips25_sap3/net1275
+ sg13g2_dlygate4sd3_1
XFILLER_33_56 VPWR VGND sg13g2_fill_1
XFILLER_20_470 VPWR VGND sg13g2_fill_1
XFILLER_4_625 VPWR VGND sg13g2_fill_2
XFILLER_3_102 VPWR VGND sg13g2_decap_4
XFILLER_3_168 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3600_ heichips25_sap3/_1173_ heichips25_sap3/_1172_ heichips25_sap3/_1056_
+ heichips25_sap3/net94 heichips25_sap3__3971_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3531_ heichips25_sap3/_1122_ heichips25_sap3/net96 heichips25_sap3/_1019_
+ VPWR VGND sg13g2_nand2_1
XFILLER_3_179 VPWR VGND sg13g2_fill_1
XFILLER_0_831 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3462_ heichips25_sap3/_0935_ heichips25_sap3/net98 heichips25_sap3/_1065_
+ VPWR VGND heichips25_sap3/_0934_ sg13g2_nand3b_1
Xheichips25_sap3__2413_ heichips25_sap3/_1734_ heichips25_sap3/_1824_ heichips25_sap3/_1828_
+ heichips25_sap3/_1829_ heichips25_sap3/_1830_ VPWR VGND sg13g2_and4_1
Xheichips25_sap3__3393_ VGND VPWR heichips25_sap3/_0976_ heichips25_sap3/_0991_ heichips25_sap3/_1001_
+ heichips25_sap3/_0999_ sg13g2_a21oi_1
Xheichips25_sap3__2344_ VGND VPWR heichips25_sap3/net224 heichips25_sap3/_1709_ heichips25_sap3/_1765_
+ heichips25_sap3/net220 sg13g2_a21oi_1
XFILLER_28_592 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2275_ heichips25_sap3/_1696_ heichips25_sap3/_1541_ heichips25_sap3/_1627_
+ VPWR VGND sg13g2_nand2_1
XFILLER_16_754 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__4014_ heichips25_sap3/net438 VGND VPWR heichips25_sap3/_0155_ heichips25_sap3__4014_/Q
+ heichips25_sap3__4014_/CLK sg13g2_dfrbpq_1
XFILLER_43_573 VPWR VGND sg13g2_fill_2
XFILLER_31_724 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2942__568 VPWR VGND net567 sg13g2_tiehi
XFILLER_30_267 VPWR VGND sg13g2_decap_8
XFILLER_7_430 VPWR VGND sg13g2_fill_2
XFILLER_8_986 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3729_ heichips25_sap3/_1246_ heichips25_sap3/_0291_ heichips25_sap3/_1245_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_can_lehmann_fsm__2950_ net535 VGND VPWR heichips25_can_lehmann_fsm/net1061
+ heichips25_can_lehmann_fsm__2950_/Q clknet_leaf_5_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2881_ net733 VGND VPWR heichips25_can_lehmann_fsm/net1096
+ heichips25_can_lehmann_fsm__2881_/Q clknet_leaf_9_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1901_ heichips25_can_lehmann_fsm/_1090_ VPWR heichips25_can_lehmann_fsm/_1214_
+ VGND heichips25_can_lehmann_fsm/net219 heichips25_can_lehmann_fsm/_1213_ sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__1832_ VGND VPWR heichips25_can_lehmann_fsm/net343 net4
+ heichips25_can_lehmann_fsm/_1148_ heichips25_can_lehmann_fsm__3044_/Q sg13g2_a21oi_1
XFILLER_0_1013 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1763_ heichips25_can_lehmann_fsm/_1081_ heichips25_can_lehmann_fsm/_1032_
+ heichips25_can_lehmann_fsm/net344 heichips25_can_lehmann_fsm/_1031_ heichips25_can_lehmann_fsm/net351
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm_hold1007 heichips25_can_lehmann_fsm__2845_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1006 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1029 heichips25_can_lehmann_fsm/_0180_ VPWR VGND heichips25_can_lehmann_fsm/net1028
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__1694_ heichips25_can_lehmann_fsm/_1018_ heichips25_can_lehmann_fsm/net296
+ heichips25_can_lehmann_fsm__2896_/Q heichips25_can_lehmann_fsm/net317 heichips25_can_lehmann_fsm__2992_/Q
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm_hold1018 heichips25_can_lehmann_fsm__2961_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1017 sg13g2_dlygate4sd3_1
XFILLER_22_713 VPWR VGND sg13g2_fill_2
XFILLER_21_234 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2315_ VGND VPWR heichips25_can_lehmann_fsm/_0607_ heichips25_can_lehmann_fsm/net1169
+ heichips25_can_lehmann_fsm/_0058_ heichips25_can_lehmann_fsm/_0622_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2246_ heichips25_can_lehmann_fsm/net170 heichips25_can_lehmann_fsm/_0566_
+ heichips25_can_lehmann_fsm/_0567_ VPWR VGND sg13g2_nor2_1
Xheichips25_can_lehmann_fsm__2177_ VPWR VGND heichips25_can_lehmann_fsm/net164 heichips25_can_lehmann_fsm/_0512_
+ heichips25_can_lehmann_fsm/_0511_ net14 heichips25_can_lehmann_fsm/_0513_ heichips25_can_lehmann_fsm/_0499_
+ sg13g2_a221oi_1
XFILLER_0_105 VPWR VGND sg13g2_decap_8
Xheichips25_sap3_fanout440 heichips25_sap3/net442 heichips25_sap3/net440 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout451 heichips25_sap3/net454 heichips25_sap3/net451 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout462 heichips25_sap3/net463 heichips25_sap3/net462 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3__2060_ heichips25_sap3/_1481_ heichips25_sap3/net234 heichips25_sap3/_1480_
+ VPWR VGND sg13g2_nand2_1
XFILLER_44_88 VPWR VGND sg13g2_fill_2
Xheichips25_sap3_hold1073 heichips25_sap3/_1356_ VPWR VGND heichips25_sap3/net1072
+ sg13g2_dlygate4sd3_1
XFILLER_12_223 VPWR VGND sg13g2_decap_8
XFILLER_9_739 VPWR VGND sg13g2_fill_1
XFILLER_12_278 VPWR VGND sg13g2_decap_8
XFILLER_21_790 VPWR VGND sg13g2_fill_1
XFILLER_5_901 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2962_ heichips25_sap3/_0599_ VPWR heichips25_sap3/_0600_ VGND heichips25_sap3/_1869_
+ heichips25_sap3/_0587_ sg13g2_o21ai_1
XFILLER_5_967 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2893_ heichips25_sap3/_0529_ VPWR heichips25_sap3/_0534_ VGND heichips25_sap3/_0532_
+ heichips25_sap3/_0533_ sg13g2_o21ai_1
XFILLER_39_109 VPWR VGND sg13g2_decap_8
XFILLER_0_672 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3514_ heichips25_sap3/_1108_ heichips25_sap3/_1096_ heichips25_sap3/_0328_
+ heichips25_sap3/_0882_ heichips25_sap3/net45 VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3445_ VGND VPWR heichips25_sap3/_1044_ heichips25_sap3/_1047_ heichips25_sap3/_1051_
+ heichips25_sap3/_1050_ sg13g2_a21oi_1
XFILLER_10_8 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2913__670 VPWR VGND net669 sg13g2_tiehi
XFILLER_36_827 VPWR VGND sg13g2_fill_1
Xclkbuf_2_3__f_clk clknet_2_3__leaf_clk clknet_0_clk VPWR VGND sg13g2_buf_16
Xheichips25_sap3__3376_ heichips25_sap3/_0076_ heichips25_sap3/_0975_ heichips25_sap3/_0982_
+ heichips25_sap3/net55 heichips25_sap3/_1400_ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2327_ heichips25_sap3/_1748_ heichips25_sap3/net73 heichips25_sap3__4002_/Q
+ heichips25_sap3/net83 heichips25_sap3__3962_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2258_ heichips25_sap3/_1679_ heichips25_sap3/net247 heichips25_sap3/_1460_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__2189_ heichips25_sap3/_1599_ heichips25_sap3/_1600_ heichips25_sap3/_1601_
+ heichips25_sap3/_1609_ heichips25_sap3/_1610_ VPWR VGND sg13g2_nor4_1
Xheichips25_can_lehmann_fsm__2100_ VGND VPWR heichips25_can_lehmann_fsm/_0438_ heichips25_can_lehmann_fsm/_0439_
+ heichips25_can_lehmann_fsm/_0025_ heichips25_can_lehmann_fsm/_0440_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2031_ heichips25_can_lehmann_fsm__2782_/Q heichips25_can_lehmann_fsm/_0312_
+ heichips25_can_lehmann_fsm/_0382_ VPWR VGND sg13g2_nor2_1
XFILLER_39_654 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2933_ net603 VGND VPWR heichips25_can_lehmann_fsm/_0158_
+ heichips25_can_lehmann_fsm__2933_/Q clknet_leaf_15_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2864_ net767 VGND VPWR heichips25_can_lehmann_fsm/net1086
+ heichips25_can_lehmann_fsm__2864_/Q clknet_leaf_8_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2795_ net616 VGND VPWR heichips25_can_lehmann_fsm/_0020_
+ heichips25_can_lehmann_fsm__2795_/Q clknet_leaf_2_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1815_ heichips25_can_lehmann_fsm/_1128_ heichips25_can_lehmann_fsm/_1124_
+ heichips25_can_lehmann_fsm/_1129_ heichips25_can_lehmann_fsm/_1131_ VPWR VGND sg13g2_a21o_1
Xheichips25_can_lehmann_fsm__1746_ heichips25_can_lehmann_fsm__2784_/Q heichips25_can_lehmann_fsm__2783_/Q
+ heichips25_can_lehmann_fsm__2782_/Q heichips25_can_lehmann_fsm__2781_/Q heichips25_can_lehmann_fsm/_1066_
+ VPWR VGND sg13g2_nor4_1
XFILLER_14_69 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1677_ heichips25_can_lehmann_fsm/net350 heichips25_can_lehmann_fsm/net351
+ heichips25_can_lehmann_fsm/net354 heichips25_can_lehmann_fsm/_1001_ VPWR VGND sg13g2_or3_1
Xheichips25_can_lehmann_fsm__2229_ VGND VPWR heichips25_can_lehmann_fsm/net162 heichips25_can_lehmann_fsm/_0552_
+ heichips25_can_lehmann_fsm/_0041_ heichips25_can_lehmann_fsm/_0553_ sg13g2_a21oi_1
XFILLER_30_79 VPWR VGND sg13g2_decap_8
XFILLER_2_937 VPWR VGND sg13g2_decap_8
XFILLER_17_304 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3230_ heichips25_sap3/_0717_ heichips25_sap3/net150 heichips25_sap3__4020_/Q
+ heichips25_sap3/_0843_ VPWR VGND sg13g2_nand3_1
XFILLER_29_131 VPWR VGND sg13g2_fill_1
XFILLER_17_315 VPWR VGND sg13g2_fill_2
XFILLER_18_849 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3161_ heichips25_sap3/_0769_ heichips25_sap3/_0773_ heichips25_sap3/_0774_
+ VPWR VGND sg13g2_and2_1
Xheichips25_sap3__2112_ heichips25_sap3/_1474_ heichips25_sap3/_1517_ heichips25_sap3/_1530_
+ heichips25_sap3/_1531_ heichips25_sap3/_1533_ VPWR VGND sg13g2_nor4_1
Xheichips25_sap3__3092_ heichips25_sap3/_0705_ heichips25_sap3/net235 heichips25_sap3/net222
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3_fanout292 heichips25_sap3/_1266_ heichips25_sap3/net292 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3__2043_ heichips25_sap3/_1464_ heichips25_sap3/net253 heichips25_sap3/net252
+ VPWR VGND sg13g2_nand2b_1
Xheichips25_sap3_fanout270 heichips25_sap3/net271 heichips25_sap3/net270 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout281 heichips25_sap3__3903_/Q heichips25_sap3/net281 VPWR VGND
+ sg13g2_buf_1
XFILLER_9_569 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3994_ heichips25_sap3/net444 VGND VPWR heichips25_sap3/_0135_ heichips25_sap3__3994_/Q
+ heichips25_sap3__4024_/CLK sg13g2_dfrbpq_1
Xheichips25_sap3__2945_ heichips25_sap3/net69 heichips25_sap3/net277 heichips25_sap3/_0583_
+ heichips25_sap3/_0046_ VPWR VGND sg13g2_a21o_1
XFILLER_4_285 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2876_ heichips25_sap3/net69 heichips25_sap3/net283 heichips25_sap3/_0517_
+ heichips25_sap3/_0043_ VPWR VGND sg13g2_a21o_1
XFILLER_0_480 VPWR VGND sg13g2_decap_4
XFILLER_0_491 VPWR VGND sg13g2_decap_8
XFILLER_49_996 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3428_ heichips25_sap3/_1034_ heichips25_sap3/net136 heichips25_sap3__3970_/Q
+ heichips25_sap3/_0768_ heichips25_sap3__3978_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_36_624 VPWR VGND sg13g2_fill_2
XFILLER_35_112 VPWR VGND sg13g2_fill_2
XFILLER_35_101 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2846__804 VPWR VGND net803 sg13g2_tiehi
XFILLER_24_819 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3359_ heichips25_sap3/_0943_ heichips25_sap3/_0965_ heichips25_sap3/_0968_
+ VPWR VGND sg13g2_and2_1
Xheichips25_can_lehmann_fsm__2580_ heichips25_can_lehmann_fsm/net478 VPWR heichips25_can_lehmann_fsm/_0756_
+ VGND heichips25_can_lehmann_fsm__2964_/Q heichips25_can_lehmann_fsm/net369 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__1600_ VPWR heichips25_can_lehmann_fsm/_0924_ heichips25_can_lehmann_fsm/net937
+ VGND sg13g2_inv_1
XFILLER_23_307 VPWR VGND sg13g2_fill_1
XFILLER_23_318 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1531_ VPWR heichips25_can_lehmann_fsm/_0855_ heichips25_can_lehmann_fsm/net1051
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__3063_ net686 VGND VPWR heichips25_can_lehmann_fsm/net1214
+ heichips25_can_lehmann_fsm__3063_/Q clknet_leaf_0_clk sg13g2_dfrbpq_1
X_26__512 VPWR VGND net511 sg13g2_tielo
Xfanout504 net506 net504 VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm__2014_ heichips25_can_lehmann_fsm/net321 VPWR heichips25_can_lehmann_fsm/_0368_
+ VGND heichips25_can_lehmann_fsm/net1240 heichips25_can_lehmann_fsm/net178 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2916_ net663 VGND VPWR heichips25_can_lehmann_fsm/net862
+ heichips25_can_lehmann_fsm__2916_/Q clknet_leaf_17_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2847_ net801 VGND VPWR heichips25_can_lehmann_fsm/_0072_
+ heichips25_can_lehmann_fsm__2847_/Q clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_41_148 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2778_ net650 VGND VPWR heichips25_can_lehmann_fsm/net1263
+ heichips25_can_lehmann_fsm__2778_/Q clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_23_830 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1729_ heichips25_can_lehmann_fsm__2829_/Q heichips25_can_lehmann_fsm__2828_/Q
+ heichips25_can_lehmann_fsm/_1050_ VPWR VGND sg13g2_nor2_1
XFILLER_22_362 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2897__702 VPWR VGND net701 sg13g2_tiehi
XFILLER_41_34 VPWR VGND sg13g2_decap_8
XFILLER_6_517 VPWR VGND sg13g2_decap_8
XFILLER_41_78 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2730_ heichips25_sap3/_0374_ heichips25_sap3/_0375_ heichips25_sap3/_0376_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__2661_ heichips25_sap3/_0323_ heichips25_sap3/_0325_ heichips25_sap3/_0005_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__2592_ heichips25_sap3/_0265_ heichips25_sap3/net71 heichips25_sap3__3981_/Q
+ heichips25_sap3/net218 heichips25_sap3__4013_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_17_123 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3213_ heichips25_sap3/_0826_ heichips25_sap3/net105 heichips25_sap3__3947_/Q
+ heichips25_sap3/net128 heichips25_sap3__3939_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3144_ heichips25_sap3/net152 heichips25_sap3/net150 heichips25_sap3/_0757_
+ VPWR VGND sg13g2_and2_1
XFILLER_9_300 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3075_ heichips25_sap3/_1548_ heichips25_sap3/_1497_ heichips25_sap3/_1518_
+ heichips25_sap3/_0688_ VPWR VGND sg13g2_a21o_1
XFILLER_13_351 VPWR VGND sg13g2_fill_2
XFILLER_41_693 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2026_ heichips25_sap3/net257 heichips25_sap3/_1446_ heichips25_sap3/_1447_
+ VPWR VGND sg13g2_nor2_1
XFILLER_9_322 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2798__611 VPWR VGND net610 sg13g2_tiehi
Xheichips25_can_lehmann_fsm_hold1190 heichips25_can_lehmann_fsm/_0618_ VPWR VGND heichips25_can_lehmann_fsm/net1189
+ sg13g2_dlygate4sd3_1
XFILLER_9_377 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3977_ heichips25_sap3/net459 VGND VPWR heichips25_sap3/_0118_ heichips25_sap3__3977_/Q
+ heichips25_sap3__3993_/CLK sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm_fanout409 heichips25_can_lehmann_fsm/net411 heichips25_can_lehmann_fsm/net409
+ VPWR VGND sg13g2_buf_1
Xheichips25_sap3__2928_ heichips25_sap3/_0567_ heichips25_sap3/_0449_ heichips25_sap3/_0349_
+ heichips25_sap3/_0416_ heichips25_sap3/net274 VPWR VGND sg13g2_a22oi_1
XFILLER_49_4 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2859_ heichips25_sap3/_1367_ heichips25_sap3/_1619_ heichips25_sap3/_1714_
+ heichips25_sap3/_0501_ VPWR VGND sg13g2_nor3_1
XFILLER_49_793 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2701_ VGND VPWR heichips25_can_lehmann_fsm/_0870_ heichips25_can_lehmann_fsm/net424
+ heichips25_can_lehmann_fsm/_0250_ heichips25_can_lehmann_fsm/_0816_ sg13g2_a21oi_1
XFILLER_36_487 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2632_ heichips25_can_lehmann_fsm/net479 VPWR heichips25_can_lehmann_fsm/_0782_
+ VGND heichips25_can_lehmann_fsm__2990_/Q heichips25_can_lehmann_fsm/net361 sg13g2_o21ai_1
XFILLER_17_690 VPWR VGND sg13g2_fill_2
XFILLER_23_115 VPWR VGND sg13g2_fill_1
XFILLER_24_649 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2563_ VGND VPWR heichips25_can_lehmann_fsm/_0907_ heichips25_can_lehmann_fsm/net427
+ heichips25_can_lehmann_fsm/_0181_ heichips25_can_lehmann_fsm/_0747_ sg13g2_a21oi_1
Xclkbuf_4_4_0_heichips25_sap3\_sap_3_inst.alu_inst.clk clknet_0_heichips25_sap3\/sap_3_inst.alu_inst.clk
+ clknet_4_4_0_heichips25_sap3\/sap_3_inst.alu_inst.clk VPWR VGND sg13g2_buf_8
Xheichips25_can_lehmann_fsm__2494_ heichips25_can_lehmann_fsm/net467 VPWR heichips25_can_lehmann_fsm/_0713_
+ VGND heichips25_can_lehmann_fsm/net962 heichips25_can_lehmann_fsm/net390 sg13g2_o21ai_1
XFILLER_11_48 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__3046_ net662 VGND VPWR heichips25_can_lehmann_fsm/_0271_
+ heichips25_can_lehmann_fsm__3046_/Q clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_47_719 VPWR VGND sg13g2_fill_1
XFILLER_36_67 VPWR VGND sg13g2_fill_2
XFILLER_15_627 VPWR VGND sg13g2_fill_1
XFILLER_11_833 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3900_ heichips25_sap3/net447 VGND VPWR heichips25_sap3/_0041_ heichips25_sap3__3900_/Q
+ heichips25_sap3__4021_/CLK sg13g2_dfrbpq_1
XFILLER_7_837 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3831_ heichips25_sap3/_1336_ heichips25_sap3/_1278_ heichips25_sap3__4010_/Q
+ heichips25_sap3/_1274_ heichips25_sap3__3946_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3762_ heichips25_sap3__4043_/Q heichips25_sap3__4042_/Q heichips25_sap3/_1271_
+ heichips25_sap3/_1274_ VPWR VGND sg13g2_nor3_1
XFILLER_7_0 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2938__584 VPWR VGND net583 sg13g2_tiehi
Xheichips25_sap3__2713_ VGND VPWR heichips25_sap3/_0359_ heichips25_sap3__3918_/Q
+ heichips25_sap3/net282 sg13g2_or2_1
Xheichips25_sap3__3693_ heichips25_sap3/_0149_ heichips25_sap3/_1140_ heichips25_sap3/_1228_
+ heichips25_sap3/_0755_ heichips25_sap3/_1406_ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2644_ VGND VPWR heichips25_sap3/_1576_ heichips25_sap3/_0307_ heichips25_sap3/_0311_
+ heichips25_sap3/_0310_ sg13g2_a21oi_1
Xheichips25_sap3__2575_ heichips25_sap3/_1695_ heichips25_sap3/_1712_ heichips25_sap3__3957_/Q
+ heichips25_sap3/_0248_ VPWR VGND heichips25_sap3/_1731_ sg13g2_nand4_1
XFILLER_46_785 VPWR VGND sg13g2_fill_1
XFILLER_45_284 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3127_ heichips25_sap3/_1485_ VPWR heichips25_sap3/_0740_ VGND heichips25_sap3/_1664_
+ heichips25_sap3/_0669_ sg13g2_o21ai_1
XFILLER_21_608 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3058_ heichips25_sap3/_0671_ heichips25_sap3/_0670_ heichips25_sap3/_0641_
+ heichips25_sap3/_0668_ heichips25_sap3/net225 VPWR VGND sg13g2_a22oi_1
XFILLER_20_129 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2009_ heichips25_sap3/_1432_ heichips25_sap3/net1130 heichips25_sap3/net835
+ VPWR VGND sg13g2_nand2_1
XFILLER_9_141 VPWR VGND sg13g2_fill_1
XFILLER_9_163 VPWR VGND sg13g2_fill_1
XFILLER_9_174 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm_fanout206 heichips25_can_lehmann_fsm/net209 heichips25_can_lehmann_fsm/net206
+ VPWR VGND sg13g2_buf_1
XFILLER_49_590 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1994_ VPWR VGND heichips25_can_lehmann_fsm/net194 heichips25_can_lehmann_fsm/_0350_
+ heichips25_can_lehmann_fsm/_0349_ heichips25_can_lehmann_fsm/_0346_ heichips25_can_lehmann_fsm/_0009_
+ heichips25_can_lehmann_fsm/_0348_ sg13g2_a221oi_1
XFILLER_37_796 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2615_ VGND VPWR heichips25_can_lehmann_fsm/_0894_ heichips25_can_lehmann_fsm/net413
+ heichips25_can_lehmann_fsm/_0207_ heichips25_can_lehmann_fsm/_0773_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2546_ heichips25_can_lehmann_fsm/net467 VPWR heichips25_can_lehmann_fsm/_0739_
+ VGND heichips25_can_lehmann_fsm/net1037 heichips25_can_lehmann_fsm/net392 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__3059__719 VPWR VGND net718 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2477_ VGND VPWR heichips25_can_lehmann_fsm/_0928_ heichips25_can_lehmann_fsm/net374
+ heichips25_can_lehmann_fsm/_0138_ heichips25_can_lehmann_fsm/_0704_ sg13g2_a21oi_1
XFILLER_0_7 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__3029_ net645 VGND VPWR heichips25_can_lehmann_fsm/_0254_
+ heichips25_can_lehmann_fsm__3029_/Q clknet_leaf_15_clk sg13g2_dfrbpq_1
Xheichips25_sap3__2360_ heichips25_sap3/_1780_ VPWR heichips25_sap3/_1781_ VGND heichips25_sap3/_1621_
+ heichips25_sap3/_1773_ sg13g2_o21ai_1
XFILLER_43_700 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2291_ VGND VPWR heichips25_sap3/_1707_ heichips25_sap3/_1708_ heichips25_sap3/_1712_
+ heichips25_sap3/_1711_ sg13g2_a21oi_1
XFILLER_27_262 VPWR VGND sg13g2_decap_8
XFILLER_28_785 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__4030_ heichips25_sap3/net461 VGND VPWR heichips25_sap3/_0171_ heichips25_sap3__4030_/Q
+ clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_43_722 VPWR VGND sg13g2_fill_1
XFILLER_42_210 VPWR VGND sg13g2_decap_8
XFILLER_27_295 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm_hold851 heichips25_can_lehmann_fsm/_0248_ VPWR VGND heichips25_can_lehmann_fsm/net850
+ sg13g2_dlygate4sd3_1
Xclkbuf_leaf_22_clk clknet_2_0__leaf_clk clknet_leaf_22_clk VPWR VGND sg13g2_buf_8
Xheichips25_can_lehmann_fsm_hold862 heichips25_can_lehmann_fsm__2915_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net861 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold884 heichips25_can_lehmann_fsm__2865_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net883 sg13g2_dlygate4sd3_1
XFILLER_11_663 VPWR VGND sg13g2_decap_8
XFILLER_11_674 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm_hold895 heichips25_can_lehmann_fsm/_0149_ VPWR VGND heichips25_can_lehmann_fsm/net894
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold873 heichips25_can_lehmann_fsm__2979_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net872 sg13g2_dlygate4sd3_1
XFILLER_6_122 VPWR VGND sg13g2_decap_4
XFILLER_6_111 VPWR VGND sg13g2_fill_2
XFILLER_10_162 VPWR VGND sg13g2_decap_8
XFILLER_10_173 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3814_ VGND VPWR heichips25_sap3__3992_/Q heichips25_sap3/net293
+ heichips25_sap3/_1321_ heichips25_sap3/net291 sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2953__813 VPWR VGND net812 sg13g2_tiehi
Xheichips25_sap3__3745_ heichips25_sap3/_1257_ heichips25_sap3__4042_/Q heichips25_sap3__4043_/Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_40_8 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3676_ VGND VPWR heichips25_sap3/_1216_ heichips25_sap3/_1217_ heichips25_sap3/_1219_
+ heichips25_sap3/_1218_ sg13g2_a21oi_1
Xheichips25_sap3__2627_ heichips25_sap3/_1455_ heichips25_sap3/_0294_ heichips25_sap3__4069_/A
+ VPWR VGND sg13g2_nor2_1
XFILLER_38_549 VPWR VGND sg13g2_fill_1
X_13_ uo_out_fsm\[7\] net524 net507 net42 VPWR VGND sg13g2_mux2_1
Xheichips25_sap3__2558_ heichips25_sap3/_0233_ heichips25_sap3/_1788_ heichips25_sap3__3891_/Q
+ heichips25_sap3/_1770_ net6 VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2489_ heichips25_sap3/_1902_ heichips25_sap3/net74 heichips25_sap3__3996_/Q
+ heichips25_sap3/net78 heichips25_sap3__4012_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_15_980 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2400_ heichips25_can_lehmann_fsm/net471 VPWR heichips25_can_lehmann_fsm/_0666_
+ VGND heichips25_can_lehmann_fsm__2875_/Q heichips25_can_lehmann_fsm/net402 sg13g2_o21ai_1
Xclkbuf_leaf_13_clk clknet_2_0__leaf_clk clknet_leaf_13_clk VPWR VGND sg13g2_buf_8
Xheichips25_can_lehmann_fsm__2331_ VGND VPWR heichips25_can_lehmann_fsm/_0969_ heichips25_can_lehmann_fsm/net403
+ heichips25_can_lehmann_fsm/_0065_ heichips25_can_lehmann_fsm/_0631_ sg13g2_a21oi_1
XFILLER_30_983 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2262_ heichips25_can_lehmann_fsm/net173 heichips25_can_lehmann_fsm/_0579_
+ heichips25_can_lehmann_fsm/_0580_ VPWR VGND sg13g2_nor2_1
Xheichips25_can_lehmann_fsm__2193_ VPWR VGND net17 heichips25_can_lehmann_fsm/_0497_
+ heichips25_can_lehmann_fsm/_0499_ heichips25_can_lehmann_fsm/net1113 heichips25_can_lehmann_fsm/_0526_
+ heichips25_can_lehmann_fsm/net175 sg13g2_a221oi_1
Xheichips25_can_lehmann_fsm__2854__788 VPWR VGND net787 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__1977_ heichips25_can_lehmann_fsm/_0336_ heichips25_can_lehmann_fsm/net187
+ heichips25_can_lehmann_fsm/_0335_ heichips25_can_lehmann_fsm/net199 heichips25_can_lehmann_fsm__2781_/Q
+ VPWR VGND sg13g2_a22oi_1
XFILLER_37_571 VPWR VGND sg13g2_fill_2
XFILLER_25_711 VPWR VGND sg13g2_fill_1
XFILLER_24_221 VPWR VGND sg13g2_decap_8
XFILLER_24_243 VPWR VGND sg13g2_fill_2
XFILLER_12_405 VPWR VGND sg13g2_decap_8
Xheichips25_sap3_hold1277 heichips25_sap3/_0007_ VPWR VGND heichips25_sap3/net1276
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__2529_ VGND VPWR heichips25_can_lehmann_fsm/_0915_ heichips25_can_lehmann_fsm/net370
+ heichips25_can_lehmann_fsm/_0164_ heichips25_can_lehmann_fsm/_0730_ sg13g2_a21oi_1
XFILLER_3_147 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3530_ heichips25_sap3/_0093_ heichips25_sap3/_1120_ heichips25_sap3/_1121_
+ heichips25_sap3/net107 heichips25_sap3/_1410_ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3461_ VGND VPWR heichips25_sap3/net122 heichips25_sap3/_0914_ heichips25_sap3/_1064_
+ net44 sg13g2_a21oi_1
XFILLER_47_346 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2412_ heichips25_sap3/_1829_ heichips25_sap3/_1745_ heichips25_sap3__4000_/Q
+ heichips25_sap3/_1743_ heichips25_sap3__4016_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3392_ heichips25_sap3/_0857_ heichips25_sap3/_0951_ heichips25_sap3/net54
+ heichips25_sap3/_1000_ VPWR VGND heichips25_sap3/_0998_ sg13g2_nand4_1
Xheichips25_sap3__2343_ heichips25_sap3/_1760_ heichips25_sap3/_1761_ heichips25_sap3/_1758_
+ heichips25_sap3/_1764_ VPWR VGND heichips25_sap3/_1763_ sg13g2_nand4_1
Xheichips25_sap3__2274_ heichips25_sap3/_1680_ heichips25_sap3/_1693_ heichips25_sap3/_1695_
+ VPWR VGND sg13g2_nor2_1
XFILLER_15_221 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__4013_ heichips25_sap3/net433 VGND VPWR heichips25_sap3/_0154_ heichips25_sap3__4013_/Q
+ heichips25_sap3__4013_/CLK sg13g2_dfrbpq_1
XFILLER_15_265 VPWR VGND sg13g2_decap_8
X_13__525 VPWR VGND net524 sg13g2_tielo
XFILLER_31_747 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__1989_ VPWR heichips25_sap3/_1415_ heichips25_sap3__4001_/Q VGND
+ sg13g2_inv_1
Xheichips25_sap3__3728_ heichips25_sap3/_1245_ heichips25_sap3/_1360_ heichips25_sap3/net832
+ VPWR VGND sg13g2_nand2_1
XFILLER_2_180 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_2_clk clknet_2_1__leaf_clk clknet_leaf_2_clk VPWR VGND sg13g2_buf_8
XFILLER_38_302 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1900_ VGND VPWR heichips25_can_lehmann_fsm/_0946_ heichips25_can_lehmann_fsm/net302
+ heichips25_can_lehmann_fsm/_1213_ heichips25_can_lehmann_fsm/_1212_ sg13g2_a21oi_1
Xheichips25_sap3__3659_ heichips25_sap3/_0138_ heichips25_sap3/_0929_ heichips25_sap3/_1205_
+ heichips25_sap3/net112 heichips25_sap3/_1377_ VPWR VGND sg13g2_a22oi_1
XFILLER_39_858 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2880_ net735 VGND VPWR heichips25_can_lehmann_fsm/net1001
+ heichips25_can_lehmann_fsm__2880_/Q clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_17_2 VPWR VGND sg13g2_fill_1
XFILLER_38_357 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1831_ heichips25_can_lehmann_fsm__3044_/Q heichips25_can_lehmann_fsm/_1145_
+ heichips25_can_lehmann_fsm__3045_/Q heichips25_can_lehmann_fsm/_1147_ VPWR VGND
+ heichips25_can_lehmann_fsm/_1146_ sg13g2_nand4_1
Xheichips25_can_lehmann_fsm__1762_ heichips25_can_lehmann_fsm/_1080_ heichips25_can_lehmann_fsm__2791_/Q
+ heichips25_can_lehmann_fsm/_1037_ VPWR VGND sg13g2_nand2_1
XFILLER_0_72 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm_hold1008 heichips25_can_lehmann_fsm/_0070_ VPWR VGND heichips25_can_lehmann_fsm/net1007
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__1693_ heichips25_can_lehmann_fsm/_1017_ heichips25_can_lehmann_fsm/net294
+ heichips25_can_lehmann_fsm__2968_/Q heichips25_can_lehmann_fsm/net331 heichips25_can_lehmann_fsm__3040_/Q
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm_hold1019 heichips25_can_lehmann_fsm/_0186_ VPWR VGND heichips25_can_lehmann_fsm/net1018
+ sg13g2_dlygate4sd3_1
XFILLER_21_224 VPWR VGND sg13g2_fill_1
XFILLER_22_758 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2314_ heichips25_can_lehmann_fsm/net329 VPWR heichips25_can_lehmann_fsm/_0622_
+ VGND heichips25_can_lehmann_fsm/net883 heichips25_can_lehmann_fsm/_0607_ sg13g2_o21ai_1
XFILLER_9_92 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2245_ heichips25_can_lehmann_fsm/_1043_ heichips25_can_lehmann_fsm/_0565_
+ heichips25_can_lehmann_fsm/_0566_ VPWR VGND sg13g2_nor2b_1
Xheichips25_can_lehmann_fsm__2176_ heichips25_can_lehmann_fsm/_0970_ heichips25_can_lehmann_fsm/_0494_
+ heichips25_can_lehmann_fsm/_0512_ VPWR VGND sg13g2_nor2_1
XFILLER_0_128 VPWR VGND sg13g2_decap_8
XFILLER_29_302 VPWR VGND sg13g2_decap_8
XFILLER_28_68 VPWR VGND sg13g2_fill_2
XFILLER_29_379 VPWR VGND sg13g2_decap_8
XFILLER_38_891 VPWR VGND sg13g2_decap_8
XFILLER_38_880 VPWR VGND sg13g2_fill_1
Xheichips25_sap3_fanout441 heichips25_sap3/net442 heichips25_sap3/net441 VPWR VGND
+ sg13g2_buf_1
XFILLER_25_530 VPWR VGND sg13g2_decap_4
XFILLER_25_552 VPWR VGND sg13g2_decap_8
Xheichips25_sap3_fanout463 _01_ heichips25_sap3/net463 VPWR VGND sg13g2_buf_1
Xheichips25_sap3_fanout452 heichips25_sap3/net453 heichips25_sap3/net452 VPWR VGND
+ sg13g2_buf_1
XFILLER_40_522 VPWR VGND sg13g2_fill_1
XFILLER_13_758 VPWR VGND sg13g2_fill_2
Xheichips25_sap3_hold1074 heichips25_sap3/_0188_ VPWR VGND heichips25_sap3/net1073
+ sg13g2_dlygate4sd3_1
XFILLER_8_239 VPWR VGND sg13g2_fill_1
XFILLER_5_924 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2961_ VPWR VGND heichips25_sap3/_0340_ heichips25_sap3/_0597_ heichips25_sap3/_0598_
+ heichips25_sap3/_0338_ heichips25_sap3/_0599_ heichips25_sap3/_0589_ sg13g2_a221oi_1
Xheichips25_sap3__2892_ heichips25_sap3/_0531_ heichips25_sap3/_0530_ heichips25_sap3/_1869_
+ heichips25_sap3/_0533_ VPWR VGND sg13g2_a21o_1
XFILLER_4_478 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3513_ heichips25_sap3/_0954_ heichips25_sap3/_1106_ heichips25_sap3/_1107_
+ VPWR VGND sg13g2_nor2b_1
Xheichips25_sap3__3444_ heichips25_sap3/_0747_ VPWR heichips25_sap3/_1050_ VGND heichips25_sap3/_1048_
+ heichips25_sap3/_1049_ sg13g2_o21ai_1
XFILLER_47_165 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3375_ heichips25_sap3/_0866_ heichips25_sap3/_0889_ heichips25_sap3/_0983_
+ heichips25_sap3/_0984_ VPWR VGND sg13g2_nor3_1
XFILLER_35_327 VPWR VGND sg13g2_decap_8
XFILLER_44_850 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2326_ VPWR VGND heichips25_sap3__3986_/Q heichips25_sap3/net90 heichips25_sap3/net75
+ heichips25_sap3__4018_/Q heichips25_sap3/_1747_ heichips25_sap3/net77 sg13g2_a221oi_1
XFILLER_18_90 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2257_ heichips25_sap3/_1470_ VPWR heichips25_sap3/_1678_ VGND heichips25_sap3/net225
+ heichips25_sap3/_1655_ sg13g2_o21ai_1
Xheichips25_sap3__2188_ heichips25_sap3/_1582_ heichips25_sap3/_1604_ heichips25_sap3/net235
+ heichips25_sap3/_1609_ VPWR VGND heichips25_sap3/_1608_ sg13g2_nand4_1
XFILLER_7_250 VPWR VGND sg13g2_decap_8
XFILLER_7_283 VPWR VGND sg13g2_fill_2
XFILLER_7_261 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2030_ heichips25_can_lehmann_fsm/_0381_ heichips25_can_lehmann_fsm/net185
+ heichips25_can_lehmann_fsm/_0380_ heichips25_can_lehmann_fsm/net198 heichips25_can_lehmann_fsm__2789_/Q
+ VPWR VGND sg13g2_a22oi_1
XFILLER_22_0 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2932_ net607 VGND VPWR heichips25_can_lehmann_fsm/_0157_
+ heichips25_can_lehmann_fsm__2932_/Q clknet_leaf_12_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2863_ net769 VGND VPWR heichips25_can_lehmann_fsm/_0088_
+ heichips25_can_lehmann_fsm__2863_/Q clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_38_154 VPWR VGND sg13g2_decap_8
XFILLER_38_143 VPWR VGND sg13g2_fill_1
XFILLER_38_132 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1814_ VGND VPWR heichips25_can_lehmann_fsm/_1124_ heichips25_can_lehmann_fsm/_1128_
+ heichips25_can_lehmann_fsm/_1130_ heichips25_can_lehmann_fsm/_1129_ sg13g2_a21oi_1
XFILLER_26_338 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2794_ net618 VGND VPWR heichips25_can_lehmann_fsm/_0019_
+ heichips25_can_lehmann_fsm__2794_/Q clknet_leaf_2_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1745_ heichips25_can_lehmann_fsm/_1065_ heichips25_can_lehmann_fsm/_1061_
+ heichips25_can_lehmann_fsm/_1064_ VPWR VGND sg13g2_nand2_1
Xheichips25_can_lehmann_fsm__1676_ heichips25_can_lehmann_fsm/net348 heichips25_can_lehmann_fsm/_0999_
+ heichips25_can_lehmann_fsm/_1000_ VPWR VGND sg13g2_nor2_1
Xclkbuf_5_14__f_heichips25_sap3\_sap_3_inst.alu_inst.clk heichips25_sap3__4024_/CLK
+ clknet_4_7_0_heichips25_sap3\/sap_3_inst.alu_inst.clk VPWR VGND sg13g2_buf_16
Xheichips25_can_lehmann_fsm__2228_ heichips25_can_lehmann_fsm/net329 VPWR heichips25_can_lehmann_fsm/_0553_
+ VGND heichips25_can_lehmann_fsm/net1221 heichips25_can_lehmann_fsm/net162 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2159_ heichips25_can_lehmann_fsm/_0493_ heichips25_can_lehmann_fsm/_0461_
+ heichips25_can_lehmann_fsm/_0494_ heichips25_can_lehmann_fsm/_0498_ VPWR VGND sg13g2_a21o_1
Xheichips25_sap3__3160_ heichips25_sap3/_0773_ heichips25_sap3/net133 heichips25_sap3__3987_/Q
+ heichips25_sap3/net134 heichips25_sap3__3963_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2111_ heichips25_sap3/net257 heichips25_sap3/_1439_ heichips25_sap3/net255
+ heichips25_sap3/_1532_ VPWR VGND sg13g2_or3_1
Xheichips25_sap3__3091_ heichips25_sap3/_0702_ VPWR heichips25_sap3/_0704_ VGND heichips25_sap3/net243
+ heichips25_sap3/_1664_ sg13g2_o21ai_1
XFILLER_26_872 VPWR VGND sg13g2_fill_1
Xheichips25_sap3_fanout293 heichips25_sap3/_1261_ heichips25_sap3/net293 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout260 heichips25_sap3__3929_/Q heichips25_sap3/net260 VPWR VGND
+ sg13g2_buf_1
XFILLER_13_522 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2042_ heichips25_sap3/net252 heichips25_sap3/net253 heichips25_sap3/_1463_
+ VPWR VGND sg13g2_nor2b_1
Xheichips25_sap3_fanout271 heichips25_sap3__3924_/Q heichips25_sap3/net271 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout282 heichips25_sap3__3902_/Q heichips25_sap3/net282 VPWR VGND
+ sg13g2_buf_1
XFILLER_9_548 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3993_ heichips25_sap3/net459 VGND VPWR heichips25_sap3/_0134_ heichips25_sap3__3993_/Q
+ heichips25_sap3__3993_/CLK sg13g2_dfrbpq_1
Xheichips25_sap3__2944_ heichips25_sap3/net69 heichips25_sap3/_0560_ heichips25_sap3/_0582_
+ heichips25_sap3/_0583_ VPWR VGND sg13g2_nor3_1
XFILLER_4_264 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2875_ VPWR VGND heichips25_sap3/_0516_ heichips25_sap3/net69 heichips25_sap3/_0515_
+ heichips25_sap3/net45 heichips25_sap3/_0517_ heichips25_sap3/net157 sg13g2_a221oi_1
XFILLER_49_942 VPWR VGND sg13g2_fill_2
XFILLER_1_982 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3427_ heichips25_sap3/_1033_ heichips25_sap3/_0772_ heichips25_sap3__3994_/Q
+ heichips25_sap3/net142 heichips25_sap3__3986_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_36_647 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3358_ heichips25_sap3/_0966_ VPWR heichips25_sap3/_0967_ VGND heichips25_sap3/net62
+ heichips25_sap3/_0944_ sg13g2_o21ai_1
Xheichips25_sap3__2309_ heichips25_sap3/_1716_ heichips25_sap3/_1728_ heichips25_sap3/_1454_
+ heichips25_sap3/_1730_ VPWR VGND heichips25_sap3/_1729_ sg13g2_nand4_1
XFILLER_16_371 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1530_ VPWR heichips25_can_lehmann_fsm/_0854_ heichips25_can_lehmann_fsm/net1043
+ VGND sg13g2_inv_1
Xheichips25_sap3__3289_ heichips25_sap3/_0901_ heichips25_sap3/_0899_ heichips25_sap3/_0858_
+ heichips25_sap3/net51 heichips25_sap3/_0859_ VPWR VGND sg13g2_a22oi_1
XFILLER_32_820 VPWR VGND sg13g2_fill_1
XFILLER_32_853 VPWR VGND sg13g2_decap_8
Xheichips25_sap3_clk_div_param_inst_hold835 heichips25_sap3_clk_div_param_inst__2_/Q
+ VPWR VGND heichips25_sap3_clk_div_param_inst__1_/A sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__3062_ net750 VGND VPWR heichips25_can_lehmann_fsm/_0287_
+ heichips25_can_lehmann_fsm__3062_/Q clknet_leaf_0_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2013_ heichips25_can_lehmann_fsm/_0366_ heichips25_can_lehmann_fsm/_0364_
+ heichips25_can_lehmann_fsm/_0365_ heichips25_can_lehmann_fsm/_0367_ VPWR VGND sg13g2_a21o_1
Xfanout505 net506 net505 VPWR VGND sg13g2_buf_1
XFILLER_39_430 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2915_ net665 VGND VPWR heichips25_can_lehmann_fsm/_0140_
+ heichips25_can_lehmann_fsm__2915_/Q clknet_leaf_17_clk sg13g2_dfrbpq_1
XFILLER_26_102 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2846_ net803 VGND VPWR heichips25_can_lehmann_fsm/_0071_
+ heichips25_can_lehmann_fsm__2846_/Q clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_26_135 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2777_ net652 VGND VPWR heichips25_can_lehmann_fsm/_0002_
+ heichips25_can_lehmann_fsm__2777_/Q clknet_leaf_14_clk sg13g2_dfrbpq_1
XFILLER_25_36 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1728_ heichips25_can_lehmann_fsm/_1046_ heichips25_can_lehmann_fsm/_1048_
+ heichips25_can_lehmann_fsm/_0973_ heichips25_can_lehmann_fsm/_1049_ VPWR VGND sg13g2_nand3_1
XFILLER_23_842 VPWR VGND sg13g2_fill_2
XFILLER_22_374 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1659_ VPWR heichips25_can_lehmann_fsm/_0983_ heichips25_can_lehmann_fsm/net348
+ VGND sg13g2_inv_1
XFILLER_10_558 VPWR VGND sg13g2_decap_8
XFILLER_1_212 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2660_ heichips25_sap3/_0325_ heichips25_sap3__4065_/Q heichips25_sap3/_1459_
+ VPWR VGND sg13g2_xnor2_1
XFILLER_1_267 VPWR VGND sg13g2_fill_2
XFILLER_49_238 VPWR VGND sg13g2_fill_2
XFILLER_1_278 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2591_ VPWR VGND heichips25_sap3__4005_/Q heichips25_sap3/net79 heichips25_sap3/net74
+ heichips25_sap3__3965_/Q heichips25_sap3/_0264_ heichips25_sap3/net83 sg13g2_a221oi_1
XFILLER_18_614 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3212_ heichips25_sap3/_0821_ heichips25_sap3/_0822_ heichips25_sap3/_0823_
+ heichips25_sap3/_0824_ heichips25_sap3/_0825_ VPWR VGND sg13g2_and4_1
Xheichips25_sap3__3143_ VPWR VGND heichips25_sap3__3995_/Q heichips25_sap3/net128
+ heichips25_sap3/net147 heichips25_sap3__4011_/Q heichips25_sap3/_0756_ heichips25_sap3/net116
+ sg13g2_a221oi_1
Xheichips25_sap3__3074_ heichips25_sap3/_1486_ heichips25_sap3/_1495_ heichips25_sap3/_1508_
+ heichips25_sap3/_0687_ VPWR VGND sg13g2_nor3_1
Xheichips25_sap3__2025_ heichips25_sap3/_1446_ heichips25_sap3/net269 heichips25_sap3/net272
+ VPWR VGND sg13g2_nand2b_1
Xheichips25_can_lehmann_fsm_hold1191 heichips25_can_lehmann_fsm/_0057_ VPWR VGND heichips25_can_lehmann_fsm/net1190
+ sg13g2_dlygate4sd3_1
XFILLER_9_367 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3976_ heichips25_sap3/net445 VGND VPWR heichips25_sap3/_0117_ heichips25_sap3__3976_/Q
+ heichips25_sap3__3993_/CLK sg13g2_dfrbpq_1
Xheichips25_sap3__2927_ heichips25_sap3/_0566_ heichips25_sap3/net278 heichips25_sap3/_0417_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__2858_ heichips25_sap3/_0500_ heichips25_sap3/_0376_ heichips25_sap3/_0378_
+ VPWR VGND sg13g2_xnor2_1
Xheichips25_sap3__2789_ heichips25_sap3/_0433_ VPWR heichips25_sap3/_0434_ VGND heichips25_sap3/_0429_
+ heichips25_sap3/_0432_ sg13g2_o21ai_1
XFILLER_37_901 VPWR VGND sg13g2_decap_4
XFILLER_49_772 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3871__816 VPWR net815 heichips25_sap3__4003_/CLK VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__2700_ heichips25_can_lehmann_fsm/net495 VPWR heichips25_can_lehmann_fsm/_0816_
+ VGND heichips25_can_lehmann_fsm__3025_/Q heichips25_can_lehmann_fsm/net424 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2631_ VGND VPWR heichips25_can_lehmann_fsm/_0890_ heichips25_can_lehmann_fsm/net395
+ heichips25_can_lehmann_fsm/_0215_ heichips25_can_lehmann_fsm/_0781_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2562_ heichips25_can_lehmann_fsm/net497 VPWR heichips25_can_lehmann_fsm/_0747_
+ VGND heichips25_can_lehmann_fsm/net1040 heichips25_can_lehmann_fsm/net427 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2493_ VGND VPWR heichips25_can_lehmann_fsm/_0924_ heichips25_can_lehmann_fsm/net356
+ heichips25_can_lehmann_fsm/_0146_ heichips25_can_lehmann_fsm/_0712_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__3045_ net678 VGND VPWR heichips25_can_lehmann_fsm/_0270_
+ heichips25_can_lehmann_fsm__3045_/Q clknet_leaf_0_clk sg13g2_dfrbpq_1
XFILLER_39_260 VPWR VGND sg13g2_decap_8
XFILLER_28_967 VPWR VGND sg13g2_decap_8
XFILLER_15_617 VPWR VGND sg13g2_decap_4
XFILLER_42_414 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2829_ net548 VGND VPWR heichips25_can_lehmann_fsm/net1166
+ heichips25_can_lehmann_fsm__2829_/Q clknet_leaf_10_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2864__768 VPWR VGND net767 sg13g2_tiehi
Xheichips25_sap3__3830_ heichips25_sap3/_1335_ heichips25_sap3/_1272_ heichips25_sap3__3978_/Q
+ heichips25_sap3/_1261_ heichips25_sap3__3994_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3761_ heichips25_sap3/_1273_ heichips25_sap3/_1272_ heichips25_sap3__3971_/Q
+ heichips25_sap3/_1270_ heichips25_sap3__4019_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2712_ heichips25_sap3/net282 heichips25_sap3__3918_/Q heichips25_sap3/_0358_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__3692_ VGND VPWR heichips25_sap3/_0888_ heichips25_sap3/_1227_ heichips25_sap3/_1228_
+ heichips25_sap3/net113 sg13g2_a21oi_1
Xheichips25_sap3__2643_ heichips25_sap3/_0310_ heichips25_sap3/_0304_ heichips25_sap3/_0308_
+ VPWR VGND sg13g2_nand2_1
XFILLER_38_709 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2574_ heichips25_sap3__3933_/Q heichips25_sap3/_1734_ heichips25_sap3/_0247_
+ VPWR VGND sg13g2_nor2_1
XFILLER_46_753 VPWR VGND sg13g2_fill_2
XFILLER_19_956 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2945__556 VPWR VGND net555 sg13g2_tiehi
Xheichips25_sap3__3126_ heichips25_sap3/_1665_ heichips25_sap3/_0646_ heichips25_sap3/_1621_
+ heichips25_sap3/_0739_ VPWR VGND heichips25_sap3/_0688_ sg13g2_nand4_1
Xheichips25_can_lehmann_fsm__3006__546 VPWR VGND net545 sg13g2_tiehi
Xheichips25_sap3__3057_ heichips25_sap3/net245 heichips25_sap3/_1515_ heichips25_sap3/_1537_
+ heichips25_sap3/_0669_ heichips25_sap3/_0670_ VPWR VGND sg13g2_nor4_1
XFILLER_14_661 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2008_ heichips25_sap3/_1431_ heichips25_sap3/net1275 heichips25_sap3/net1162
+ VPWR VGND sg13g2_nand2_1
Xheichips25_can_lehmann_fsm_fanout207 heichips25_can_lehmann_fsm/net208 heichips25_can_lehmann_fsm/net207
+ VPWR VGND sg13g2_buf_1
Xheichips25_sap3__3959_ heichips25_sap3/net459 VGND VPWR heichips25_sap3/_0100_ heichips25_sap3__3959_/Q
+ clkload29/A sg13g2_dfrbpq_1
XFILLER_47_2 VPWR VGND sg13g2_fill_1
XFILLER_3_1012 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1993_ heichips25_can_lehmann_fsm/net321 VPWR heichips25_can_lehmann_fsm/_0350_
+ VGND heichips25_can_lehmann_fsm/net1234 heichips25_can_lehmann_fsm/net177 sg13g2_o21ai_1
XFILLER_36_230 VPWR VGND sg13g2_fill_1
XFILLER_12_609 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2614_ heichips25_can_lehmann_fsm/net486 VPWR heichips25_can_lehmann_fsm/_0773_
+ VGND heichips25_can_lehmann_fsm/net1030 heichips25_can_lehmann_fsm/net413 sg13g2_o21ai_1
XFILLER_11_108 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2545_ VGND VPWR heichips25_can_lehmann_fsm/_0911_ heichips25_can_lehmann_fsm/net355
+ heichips25_can_lehmann_fsm/_0172_ heichips25_can_lehmann_fsm/_0738_ sg13g2_a21oi_1
XFILLER_20_631 VPWR VGND sg13g2_fill_1
XFILLER_20_642 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2476_ heichips25_can_lehmann_fsm/net483 VPWR heichips25_can_lehmann_fsm/_0704_
+ VGND heichips25_can_lehmann_fsm/net975 heichips25_can_lehmann_fsm/net374 sg13g2_o21ai_1
XFILLER_20_653 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__3028_ net658 VGND VPWR heichips25_can_lehmann_fsm/_0253_
+ heichips25_can_lehmann_fsm__3028_/Q clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_47_78 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2290_ heichips25_sap3/_1679_ heichips25_sap3/_1710_ heichips25_sap3/net241
+ heichips25_sap3/_1711_ VPWR VGND sg13g2_nand3_1
XFILLER_16_926 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2981__701 VPWR VGND net700 sg13g2_tiehi
XFILLER_43_712 VPWR VGND sg13g2_decap_4
XFILLER_15_414 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_hold852 heichips25_can_lehmann_fsm__2843_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net851 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold841 heichips25_can_lehmann_fsm__2851_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net840 sg13g2_dlygate4sd3_1
XFILLER_8_39 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm_hold885 heichips25_can_lehmann_fsm/_0090_ VPWR VGND heichips25_can_lehmann_fsm/net884
+ sg13g2_dlygate4sd3_1
XFILLER_7_624 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_hold863 heichips25_can_lehmann_fsm/_0141_ VPWR VGND heichips25_can_lehmann_fsm/net862
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold874 heichips25_can_lehmann_fsm/_0205_ VPWR VGND heichips25_can_lehmann_fsm/net873
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold896 heichips25_can_lehmann_fsm__2837_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net895 sg13g2_dlygate4sd3_1
Xheichips25_sap3__3813_ heichips25_sap3/_1320_ heichips25_sap3/net292 heichips25_sap3__3960_/Q
+ heichips25_sap3/_1265_ heichips25_sap3__4000_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3744_ heichips25_sap3/net836 VPWR heichips25_sap3/_0172_ VGND heichips25_sap3/_1360_
+ heichips25_sap3/_1431_ sg13g2_o21ai_1
XFILLER_2_340 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3675_ heichips25_sap3/_1218_ heichips25_sap3/net146 uio_oe_sap3\[6\]
+ VPWR VGND sg13g2_nand2b_1
XFILLER_3_885 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2626_ heichips25_sap3/_0294_ heichips25_sap3/_1784_ heichips25_sap3/_0293_
+ heichips25_sap3/net228 heichips25_sap3/net248 VPWR VGND sg13g2_a22oi_1
X_12_ uo_out_fsm\[6\] net523 net507 net41 VPWR VGND sg13g2_mux2_1
Xheichips25_sap3__2557_ VPWR VGND heichips25_sap3/_0231_ heichips25_sap3/_1654_ heichips25_sap3/_0227_
+ heichips25_sap3/_1368_ heichips25_sap3/_0232_ heichips25_sap3/net92 sg13g2_a221oi_1
XFILLER_46_550 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2488_ heichips25_sap3__3980_/Q heichips25_sap3/net76 heichips25_sap3/_1901_
+ VPWR VGND sg13g2_and2_1
XFILLER_18_274 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3109_ heichips25_sap3/net242 heichips25_sap3/_1664_ heichips25_sap3/_0295_
+ heichips25_sap3/_0722_ VPWR VGND sg13g2_nor3_1
Xheichips25_can_lehmann_fsm__2330_ heichips25_can_lehmann_fsm/net471 VPWR heichips25_can_lehmann_fsm/_0631_
+ VGND heichips25_can_lehmann_fsm/net1113 heichips25_can_lehmann_fsm/net403 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2261_ heichips25_can_lehmann_fsm/_1045_ heichips25_can_lehmann_fsm/_0578_
+ heichips25_can_lehmann_fsm/_0579_ VPWR VGND sg13g2_nor2b_1
Xheichips25_can_lehmann_fsm__2192_ heichips25_can_lehmann_fsm/net164 VPWR heichips25_can_lehmann_fsm/_0525_
+ VGND heichips25_can_lehmann_fsm/_1100_ heichips25_can_lehmann_fsm/_0524_ sg13g2_o21ai_1
Xheichips25_sap3__3877__822 VPWR net821 clkload27/A VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__1976_ heichips25_can_lehmann_fsm/_0326_ heichips25_can_lehmann_fsm/net1257
+ heichips25_can_lehmann_fsm/_0335_ VPWR VGND sg13g2_xor2_1
XFILLER_40_737 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2528_ heichips25_can_lehmann_fsm/net477 VPWR heichips25_can_lehmann_fsm/_0730_
+ VGND heichips25_can_lehmann_fsm__2938_/Q heichips25_can_lehmann_fsm/net370 sg13g2_o21ai_1
XFILLER_33_69 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2459_ VGND VPWR heichips25_can_lehmann_fsm/_0933_ heichips25_can_lehmann_fsm/net405
+ heichips25_can_lehmann_fsm/_0129_ heichips25_can_lehmann_fsm/_0695_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__3035__550 VPWR VGND net549 sg13g2_tiehi
Xheichips25_sap3__3460_ heichips25_sap3/_1060_ VPWR heichips25_sap3/_0081_ VGND heichips25_sap3/net57
+ heichips25_sap3/_1063_ sg13g2_o21ai_1
Xheichips25_sap3__2411_ heichips25_sap3/_1828_ heichips25_sap3/net72 heichips25_sap3__3976_/Q
+ heichips25_sap3/net217 heichips25_sap3__4008_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3391_ heichips25_sap3/net53 heichips25_sap3/_0857_ heichips25_sap3/_0951_
+ heichips25_sap3/_0998_ heichips25_sap3/_0999_ VPWR VGND sg13g2_and4_1
Xheichips25_sap3__2342_ heichips25_sap3/_1759_ heichips25_sap3/_1762_ heichips25_sap3/_1763_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__2273_ VPWR heichips25_sap3/_1694_ heichips25_sap3/_1693_ VGND sg13g2_inv_1
XFILLER_43_553 VPWR VGND sg13g2_fill_2
XFILLER_16_756 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__4012_ heichips25_sap3/net434 VGND VPWR heichips25_sap3/_0153_ heichips25_sap3__4012_/Q
+ heichips25_sap3__4012_/CLK sg13g2_dfrbpq_1
XFILLER_31_726 VPWR VGND sg13g2_fill_1
XFILLER_15_288 VPWR VGND sg13g2_decap_8
XFILLER_11_450 VPWR VGND sg13g2_decap_8
XFILLER_12_951 VPWR VGND sg13g2_fill_2
XFILLER_7_432 VPWR VGND sg13g2_fill_1
XFILLER_11_483 VPWR VGND sg13g2_decap_8
XFILLER_7_443 VPWR VGND sg13g2_decap_4
XFILLER_11_494 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__1988_ VPWR heichips25_sap3/_1414_ heichips25_sap3__4009_/Q VGND
+ sg13g2_inv_1
Xheichips25_sap3__3727_ VGND VPWR heichips25_sap3/net118 heichips25_sap3/_1177_ heichips25_sap3/_0167_
+ heichips25_sap3/_1244_ sg13g2_a21oi_1
XFILLER_2_170 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3658_ VPWR VGND heichips25_sap3/_1104_ heichips25_sap3/net112 heichips25_sap3/_1204_
+ heichips25_sap3/_0927_ heichips25_sap3/_1205_ heichips25_sap3/_1203_ sg13g2_a221oi_1
XFILLER_38_336 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3589_ heichips25_sap3/net136 VPWR heichips25_sap3/_1165_ VGND heichips25_sap3/_1117_
+ heichips25_sap3/_1164_ sg13g2_o21ai_1
Xheichips25_sap3__2609_ heichips25_sap3/_0280_ heichips25_sap3/_0279_ heichips25_sap3/_1528_
+ heichips25_sap3/_0278_ heichips25_sap3/_1498_ VPWR VGND sg13g2_a22oi_1
XFILLER_38_347 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__1830_ heichips25_can_lehmann_fsm/_1146_ net5 heichips25_can_lehmann_fsm/net343
+ VPWR VGND sg13g2_nand2b_1
Xheichips25_can_lehmann_fsm__1761_ uo_out_fsm\[5\] heichips25_can_lehmann_fsm/_1078_
+ heichips25_can_lehmann_fsm/_1079_ VPWR VGND sg13g2_nand2_1
XFILLER_34_553 VPWR VGND sg13g2_fill_2
XFILLER_34_542 VPWR VGND sg13g2_decap_8
XFILLER_0_84 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1692_ VGND VPWR heichips25_can_lehmann_fsm/_0951_ heichips25_can_lehmann_fsm/net300
+ heichips25_can_lehmann_fsm/_1016_ heichips25_can_lehmann_fsm/_1015_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm_hold1009 heichips25_can_lehmann_fsm__2901_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1008 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__3060__654 VPWR VGND net653 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2313_ heichips25_can_lehmann_fsm/_0620_ heichips25_can_lehmann_fsm/net1168
+ heichips25_can_lehmann_fsm/_0621_ VPWR VGND sg13g2_xor2_1
Xheichips25_can_lehmann_fsm__2244_ heichips25_can_lehmann_fsm/net1195 VPWR heichips25_can_lehmann_fsm/_0565_
+ VGND heichips25_can_lehmann_fsm__2819_/Q heichips25_can_lehmann_fsm__2818_/Q sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2175_ heichips25_can_lehmann_fsm/_1097_ heichips25_can_lehmann_fsm/net1202
+ heichips25_can_lehmann_fsm/_0511_ VPWR VGND sg13g2_xor2_1
XFILLER_29_325 VPWR VGND sg13g2_decap_8
XFILLER_29_358 VPWR VGND sg13g2_decap_8
Xheichips25_sap3_fanout442 heichips25_sap3/net446 heichips25_sap3/net442 VPWR VGND
+ sg13g2_buf_1
Xheichips25_can_lehmann_fsm__1959_ VPWR VGND heichips25_can_lehmann_fsm/net191 heichips25_can_lehmann_fsm/_0319_
+ heichips25_can_lehmann_fsm/_0320_ heichips25_can_lehmann_fsm/_0317_ heichips25_can_lehmann_fsm/_0004_
+ heichips25_can_lehmann_fsm/_0318_ sg13g2_a221oi_1
Xheichips25_sap3_hold1020 heichips25_sap3__4048_/Q VPWR VGND heichips25_sap3/net1019
+ sg13g2_dlygate4sd3_1
Xheichips25_sap3_fanout453 heichips25_sap3/net454 heichips25_sap3/net453 VPWR VGND
+ sg13g2_buf_1
XFILLER_25_575 VPWR VGND sg13g2_decap_8
XFILLER_9_719 VPWR VGND sg13g2_decap_8
XFILLER_12_258 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2960_ heichips25_sap3/_0412_ heichips25_sap3/_0410_ heichips25_sap3/_0598_
+ VPWR VGND sg13g2_xor2_1
XFILLER_20_291 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2891_ heichips25_sap3/_0530_ heichips25_sap3/_0531_ heichips25_sap3/_0532_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_can_lehmann_fsm_fanout390 heichips25_can_lehmann_fsm/net392 heichips25_can_lehmann_fsm/net390
+ VPWR VGND sg13g2_buf_1
Xheichips25_sap3__3512_ heichips25_sap3/_1106_ heichips25_sap3/net97 heichips25_sap3/_0946_
+ VPWR VGND sg13g2_nand2_1
XFILLER_47_122 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3443_ uio_oe_sap3\[7\] heichips25_sap3/_0884_ heichips25_sap3/_1049_
+ VPWR VGND sg13g2_nor2_1
XFILLER_48_678 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3374_ VGND VPWR heichips25_sap3/_0820_ heichips25_sap3/_0864_ heichips25_sap3/_0983_
+ heichips25_sap3/_0810_ sg13g2_a21oi_1
Xheichips25_sap3__2325_ heichips25_sap3/_1746_ heichips25_sap3/_1680_ heichips25_sap3/_1713_
+ heichips25_sap3/_1731_ VPWR VGND sg13g2_and3_1
XFILLER_16_520 VPWR VGND sg13g2_fill_1
XFILLER_43_361 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2256_ heichips25_sap3/_1454_ VPWR heichips25_sap3/_1677_ VGND heichips25_sap3/_1657_
+ heichips25_sap3/_1676_ sg13g2_o21ai_1
XFILLER_31_501 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2187_ heichips25_sap3/_1517_ VPWR heichips25_sap3/_1608_ VGND heichips25_sap3/_1605_
+ heichips25_sap3/_1607_ sg13g2_o21ai_1
XFILLER_31_512 VPWR VGND sg13g2_fill_1
XFILLER_31_545 VPWR VGND sg13g2_decap_8
XFILLER_4_980 VPWR VGND sg13g2_decap_8
XFILLER_38_100 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2931_ net611 VGND VPWR heichips25_can_lehmann_fsm/_0156_
+ heichips25_can_lehmann_fsm__2931_/Q clknet_leaf_12_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2862_ net771 VGND VPWR heichips25_can_lehmann_fsm/_0087_
+ heichips25_can_lehmann_fsm__2862_/Q clknet_leaf_10_clk sg13g2_dfrbpq_1
XFILLER_38_188 VPWR VGND sg13g2_fill_1
XFILLER_26_317 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1813_ heichips25_can_lehmann_fsm__2875_/Q heichips25_can_lehmann_fsm/net336
+ heichips25_can_lehmann_fsm/_1129_ VPWR VGND sg13g2_nor2_1
XFILLER_27_829 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2793_ net620 VGND VPWR heichips25_can_lehmann_fsm/net1256
+ heichips25_can_lehmann_fsm__2793_/Q clknet_leaf_4_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1744_ heichips25_can_lehmann_fsm__2780_/Q heichips25_can_lehmann_fsm__2779_/Q
+ heichips25_can_lehmann_fsm__2778_/Q heichips25_can_lehmann_fsm/_1064_ VPWR VGND
+ sg13g2_nor3_1
Xheichips25_can_lehmann_fsm__1675_ VGND VPWR heichips25_can_lehmann_fsm/_0999_ heichips25_can_lehmann_fsm/net353
+ heichips25_can_lehmann_fsm/net352 sg13g2_or2_1
XFILLER_14_38 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2227_ heichips25_can_lehmann_fsm/_0552_ heichips25_can_lehmann_fsm/net165
+ heichips25_can_lehmann_fsm/_0551_ heichips25_can_lehmann_fsm/net176 heichips25_can_lehmann_fsm/net1115
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2158_ VGND VPWR heichips25_can_lehmann_fsm/_0461_ heichips25_can_lehmann_fsm/_0493_
+ heichips25_can_lehmann_fsm/_0497_ heichips25_can_lehmann_fsm/_0494_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2089_ heichips25_can_lehmann_fsm/_0431_ heichips25_can_lehmann_fsm/_1058_
+ heichips25_can_lehmann_fsm/_0430_ VPWR VGND sg13g2_nand2_1
XFILLER_39_57 VPWR VGND sg13g2_decap_8
XFILLER_29_111 VPWR VGND sg13g2_decap_4
XFILLER_17_328 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3090_ heichips25_sap3/_0307_ VPWR heichips25_sap3/_0703_ VGND heichips25_sap3/net236
+ heichips25_sap3/_0702_ sg13g2_o21ai_1
Xheichips25_sap3__2110_ heichips25_sap3/net257 heichips25_sap3/_1439_ heichips25_sap3/net255
+ heichips25_sap3/_1531_ VPWR VGND sg13g2_nor3_1
XFILLER_13_501 VPWR VGND sg13g2_fill_2
Xheichips25_sap3_fanout250 heichips25_sap3__4066_/Q heichips25_sap3/net250 VPWR VGND
+ sg13g2_buf_1
XFILLER_41_821 VPWR VGND sg13g2_fill_1
Xheichips25_sap3_fanout272 heichips25_sap3__3923_/Q heichips25_sap3/net272 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3__2041_ heichips25_sap3/_1462_ heichips25_sap3/net247 heichips25_sap3/_1459_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3_fanout261 heichips25_sap3__3928_/Q heichips25_sap3/net261 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout283 heichips25_sap3__3902_/Q heichips25_sap3/net283 VPWR VGND
+ sg13g2_buf_1
XFILLER_41_876 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3992_ heichips25_sap3/net445 VGND VPWR heichips25_sap3/_0133_ heichips25_sap3__3992_/Q
+ clkload22/A sg13g2_dfrbpq_1
Xheichips25_sap3__2943_ VPWR VGND heichips25_sap3/_0581_ heichips25_sap3/net157 heichips25_sap3/_0580_
+ heichips25_sap3__3913_/Q heichips25_sap3/_0582_ heichips25_sap3/net203 sg13g2_a221oi_1
XFILLER_4_221 VPWR VGND sg13g2_fill_2
XFILLER_4_210 VPWR VGND sg13g2_fill_2
XFILLER_5_799 VPWR VGND sg13g2_fill_2
XFILLER_5_788 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2874_ VGND VPWR heichips25_sap3__3910_/Q heichips25_sap3/net203
+ heichips25_sap3/_0516_ heichips25_sap3/net157 sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2874__748 VPWR VGND net747 sg13g2_tiehi
XFILLER_45_1027 VPWR VGND sg13g2_fill_2
XFILLER_1_961 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3426_ heichips25_sap3/_1032_ heichips25_sap3__3962_/Q heichips25_sap3/net145
+ VPWR VGND sg13g2_nand2_1
XFILLER_36_626 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3357_ VPWR heichips25_sap3/_0966_ heichips25_sap3/_0965_ VGND sg13g2_inv_1
X_19__521 VPWR VGND net520 sg13g2_tielo
Xheichips25_sap3__2308_ heichips25_sap3/_1729_ heichips25_sap3/_1723_ heichips25_sap3/_1618_
+ heichips25_sap3/_1720_ heichips25_sap3/net272 VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3288_ heichips25_sap3/_0857_ heichips25_sap3/_0899_ heichips25_sap3/net53
+ heichips25_sap3/_0900_ VPWR VGND sg13g2_nand3_1
Xheichips25_sap3__2239_ VPWR VGND heichips25_sap3/net245 heichips25_sap3/_1577_ heichips25_sap3/_1581_
+ heichips25_sap3/net242 heichips25_sap3/_1660_ heichips25_sap3/_1559_ sg13g2_a221oi_1
XFILLER_16_361 VPWR VGND sg13g2_fill_2
XFILLER_16_383 VPWR VGND sg13g2_decap_4
XFILLER_31_331 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__3061_ net525 VGND VPWR heichips25_can_lehmann_fsm/_0286_
+ heichips25_can_lehmann_fsm__3061_/Q clknet_leaf_0_clk sg13g2_dfrbpq_1
XFILLER_6_83 VPWR VGND sg13g2_fill_2
XFILLER_6_72 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2012_ VPWR VGND heichips25_can_lehmann_fsm__2788_/Q heichips25_can_lehmann_fsm/net191
+ heichips25_can_lehmann_fsm/net188 heichips25_can_lehmann_fsm__2786_/Q heichips25_can_lehmann_fsm/_0366_
+ heichips25_can_lehmann_fsm/net197 sg13g2_a221oi_1
Xfanout506 net1 net506 VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm__2914_ net667 VGND VPWR heichips25_can_lehmann_fsm/_0139_
+ heichips25_can_lehmann_fsm__2914_/Q clknet_leaf_17_clk sg13g2_dfrbpq_1
XFILLER_27_615 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2845_ net805 VGND VPWR heichips25_can_lehmann_fsm/net1007
+ heichips25_can_lehmann_fsm__2845_/Q clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_42_629 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2776_ net654 VGND VPWR heichips25_can_lehmann_fsm/_0001_
+ heichips25_can_lehmann_fsm__2776_/Q clknet_leaf_14_clk sg13g2_dfrbpq_1
XFILLER_26_158 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1727_ heichips25_can_lehmann_fsm__2827_/Q heichips25_can_lehmann_fsm__2826_/Q
+ heichips25_can_lehmann_fsm/_1048_ VPWR VGND sg13g2_nor2_1
XFILLER_35_692 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1658_ VPWR heichips25_can_lehmann_fsm/_0982_ heichips25_can_lehmann_fsm/net1234
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__1589_ VPWR heichips25_can_lehmann_fsm/_0913_ heichips25_can_lehmann_fsm/net1025
+ VGND sg13g2_inv_1
Xheichips25_sap3__2590_ heichips25_sap3/_0263_ heichips25_sap3/net78 heichips25_sap3__4021_/Q
+ heichips25_sap3/net88 heichips25_sap3__3949_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_49_217 VPWR VGND sg13g2_decap_8
XFILLER_45_423 VPWR VGND sg13g2_fill_2
XFILLER_18_637 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3211_ heichips25_sap3/_0824_ heichips25_sap3/net133 heichips25_sap3__3995_/Q
+ heichips25_sap3/net134 heichips25_sap3__3971_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3142_ heichips25_sap3/_0755_ heichips25_sap3/_0680_ heichips25_sap3/_0717_
+ VPWR VGND sg13g2_nand2_1
XFILLER_26_692 VPWR VGND sg13g2_fill_2
XFILLER_32_128 VPWR VGND sg13g2_fill_2
XFILLER_33_629 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3073_ heichips25_sap3/net245 heichips25_sap3/_0685_ heichips25_sap3/net266
+ heichips25_sap3/_0686_ VPWR VGND sg13g2_nand3_1
Xheichips25_sap3__2024_ heichips25_sap3/net272 heichips25_sap3/net271 heichips25_sap3/_1445_
+ VPWR VGND sg13g2_nor2b_1
XFILLER_13_353 VPWR VGND sg13g2_fill_1
XFILLER_15_92 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_hold1181 heichips25_can_lehmann_fsm__2811_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1180 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1192 heichips25_can_lehmann_fsm__2826_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1191 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1170 heichips25_can_lehmann_fsm/_0621_ VPWR VGND heichips25_can_lehmann_fsm/net1169
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__2956__801 VPWR VGND net800 sg13g2_tiehi
Xheichips25_sap3__3975_ heichips25_sap3/net459 VGND VPWR heichips25_sap3/_0116_ heichips25_sap3__3975_/Q
+ clkload29/A sg13g2_dfrbpq_1
Xheichips25_sap3__2926_ heichips25_sap3/_0564_ heichips25_sap3/_0563_ heichips25_sap3/_0565_
+ VPWR VGND sg13g2_nor2b_1
Xheichips25_sap3__2857_ heichips25_sap3/_0499_ heichips25_sap3/_0449_ heichips25_sap3/_0357_
+ VPWR VGND sg13g2_nand2b_1
Xheichips25_sap3__2788_ heichips25_sap3/net228 heichips25_sap3/_1643_ heichips25_sap3/_1451_
+ heichips25_sap3/_0433_ VPWR VGND sg13g2_nand3_1
XFILLER_0_290 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3409_ heichips25_sap3/_1016_ heichips25_sap3/_0991_ heichips25_sap3/_1014_
+ VPWR VGND sg13g2_nand2_1
XFILLER_36_423 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2630_ heichips25_can_lehmann_fsm/net476 VPWR heichips25_can_lehmann_fsm/_0781_
+ VGND heichips25_can_lehmann_fsm/net1053 heichips25_can_lehmann_fsm/net395 sg13g2_o21ai_1
XFILLER_36_489 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2561_ VGND VPWR heichips25_can_lehmann_fsm/_0907_ heichips25_can_lehmann_fsm/net386
+ heichips25_can_lehmann_fsm/_0180_ heichips25_can_lehmann_fsm/_0746_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2492_ heichips25_can_lehmann_fsm/net466 VPWR heichips25_can_lehmann_fsm/_0712_
+ VGND heichips25_can_lehmann_fsm__2920_/Q heichips25_can_lehmann_fsm/net356 sg13g2_o21ai_1
XFILLER_11_17 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__3044_ net694 VGND VPWR heichips25_can_lehmann_fsm/net1230
+ heichips25_can_lehmann_fsm__3044_/Q clknet_leaf_0_clk sg13g2_dfrbpq_1
XFILLER_27_401 VPWR VGND sg13g2_fill_2
XFILLER_28_902 VPWR VGND sg13g2_fill_1
XFILLER_28_946 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2828_ net550 VGND VPWR heichips25_can_lehmann_fsm/_0053_
+ heichips25_can_lehmann_fsm__2828_/Q clknet_leaf_10_clk sg13g2_dfrbpq_1
Xclkbuf_5_15__f_heichips25_sap3\_sap_3_inst.alu_inst.clk clkload22/A clknet_4_7_0_heichips25_sap3\/sap_3_inst.alu_inst.clk
+ VPWR VGND sg13g2_buf_16
Xheichips25_can_lehmann_fsm__2759_ VGND VPWR heichips25_can_lehmann_fsm/_0855_ heichips25_can_lehmann_fsm/net419
+ heichips25_can_lehmann_fsm/_0279_ heichips25_can_lehmann_fsm/_0845_ sg13g2_a21oi_1
XFILLER_10_301 VPWR VGND sg13g2_decap_4
XFILLER_23_673 VPWR VGND sg13g2_decap_8
XFILLER_11_835 VPWR VGND sg13g2_fill_1
XFILLER_22_183 VPWR VGND sg13g2_fill_2
XFILLER_10_356 VPWR VGND sg13g2_fill_1
XFILLER_10_367 VPWR VGND sg13g2_fill_1
XFILLER_11_868 VPWR VGND sg13g2_fill_1
XFILLER_6_338 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3760_ heichips25_sap3/_1257_ heichips25_sap3/_1271_ heichips25_sap3/_1272_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__3691_ heichips25_sap3/_1227_ heichips25_sap3/_0802_ heichips25_sap3/_0867_
+ VPWR VGND sg13g2_xnor2_1
Xheichips25_sap3__2711_ heichips25_sap3/_0357_ heichips25_sap3/net282 heichips25_sap3__3918_/Q
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__2642_ heichips25_sap3/_1487_ heichips25_sap3/_1502_ heichips25_sap3/net237
+ heichips25_sap3/_0309_ VPWR VGND heichips25_sap3/_1541_ sg13g2_nand4_1
Xheichips25_sap3__2573_ heichips25_sap3/_0032_ heichips25_sap3/_0245_ heichips25_sap3/_0246_
+ VPWR VGND sg13g2_nand2_1
XFILLER_46_710 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__3012__787 VPWR VGND net786 sg13g2_tiehi
XFILLER_18_401 VPWR VGND sg13g2_fill_2
XFILLER_19_902 VPWR VGND sg13g2_decap_8
XFILLER_19_913 VPWR VGND sg13g2_fill_1
XFILLER_45_220 VPWR VGND sg13g2_decap_8
XFILLER_45_264 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3125_ VGND VPWR heichips25_sap3/_1554_ heichips25_sap3/net225 heichips25_sap3/_0738_
+ heichips25_sap3/_1536_ sg13g2_a21oi_1
Xheichips25_sap3__3056_ heichips25_sap3/_1441_ heichips25_sap3/_1495_ heichips25_sap3/_0669_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__2007_ VPWR heichips25_sap3__4062_/D heichips25_sap3/net339 VGND
+ sg13g2_inv_1
XFILLER_9_154 VPWR VGND sg13g2_decap_8
XFILLER_9_198 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm_fanout208 heichips25_can_lehmann_fsm/net209 heichips25_can_lehmann_fsm/net208
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout219 heichips25_can_lehmann_fsm/_1138_ heichips25_can_lehmann_fsm/net219
+ VPWR VGND sg13g2_buf_1
Xheichips25_sap3__3958_ heichips25_sap3/net457 VGND VPWR heichips25_sap3/_0099_ heichips25_sap3__3958_/Q
+ heichips25_sap3__3990_/CLK sg13g2_dfrbpq_1
Xheichips25_sap3__2909_ heichips25_sap3/_0408_ heichips25_sap3/_0407_ heichips25_sap3/_0549_
+ VPWR VGND sg13g2_xor2_1
Xheichips25_can_lehmann_fsm__2952__528 VPWR VGND net527 sg13g2_tiehi
Xheichips25_sap3__3889_ heichips25_sap3/net451 VGND VPWR heichips25_sap3/_0030_ heichips25_sap3__3889_/Q
+ heichips25_sap3__3921_/CLK sg13g2_dfrbpq_1
XFILLER_3_95 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1992_ heichips25_can_lehmann_fsm__2801_/Q heichips25_can_lehmann_fsm/net181
+ heichips25_can_lehmann_fsm/_0349_ VPWR VGND sg13g2_nor2_1
XFILLER_49_592 VPWR VGND sg13g2_fill_1
XFILLER_36_297 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2613_ VGND VPWR heichips25_can_lehmann_fsm/_0894_ heichips25_can_lehmann_fsm/net372
+ heichips25_can_lehmann_fsm/_0206_ heichips25_can_lehmann_fsm/_0772_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2544_ heichips25_can_lehmann_fsm/net467 VPWR heichips25_can_lehmann_fsm/_0738_
+ VGND heichips25_can_lehmann_fsm__2946_/Q heichips25_can_lehmann_fsm/net355 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2475_ VGND VPWR heichips25_can_lehmann_fsm/_0929_ heichips25_can_lehmann_fsm/net415
+ heichips25_can_lehmann_fsm/_0137_ heichips25_can_lehmann_fsm/_0703_ sg13g2_a21oi_1
XFILLER_3_319 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2900__696 VPWR VGND net695 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__3027_ net666 VGND VPWR heichips25_can_lehmann_fsm/net961
+ heichips25_can_lehmann_fsm__3027_/Q clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_47_529 VPWR VGND sg13g2_decap_4
XFILLER_27_242 VPWR VGND sg13g2_fill_2
XFILLER_15_459 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_hold853 heichips25_can_lehmann_fsm/_0069_ VPWR VGND heichips25_can_lehmann_fsm/net852
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold842 heichips25_can_lehmann_fsm/_0077_ VPWR VGND heichips25_can_lehmann_fsm/net841
+ sg13g2_dlygate4sd3_1
XFILLER_42_289 VPWR VGND sg13g2_decap_8
XFILLER_10_131 VPWR VGND sg13g2_decap_8
XFILLER_10_142 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_hold886 heichips25_can_lehmann_fsm__2967_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net885 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold875 heichips25_can_lehmann_fsm__2965_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net874 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold864 heichips25_can_lehmann_fsm__2933_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net863 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold897 heichips25_can_lehmann_fsm/_0062_ VPWR VGND heichips25_can_lehmann_fsm/net896
+ sg13g2_dlygate4sd3_1
Xheichips25_sap3__3812_ heichips25_sap3/_1319_ heichips25_sap3/_1282_ heichips25_sap3__3952_/Q
+ heichips25_sap3/_1274_ heichips25_sap3__3944_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_6_146 VPWR VGND sg13g2_decap_4
XFILLER_12_71 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3743_ heichips25_sap3/_1256_ heichips25_sap3/net835 heichips25_sap3/_1245_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__3674_ heichips25_sap3/_0889_ heichips25_sap3/_1017_ heichips25_sap3/_1217_
+ VPWR VGND sg13g2_nor2_1
XFILLER_2_396 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2625_ heichips25_sap3/_1667_ heichips25_sap3/_1775_ heichips25_sap3/_1630_
+ heichips25_sap3/_0293_ VPWR VGND heichips25_sap3/_0292_ sg13g2_nand4_1
XFILLER_26_8 VPWR VGND sg13g2_decap_8
X_11_ uo_out_fsm\[5\] uo_out_sap3\[5\] net507 net40 VPWR VGND sg13g2_mux2_1
Xheichips25_sap3__2556_ heichips25_sap3/_1734_ heichips25_sap3/_0228_ heichips25_sap3/_0229_
+ heichips25_sap3/_0230_ heichips25_sap3/_0231_ VPWR VGND sg13g2_and4_1
Xheichips25_sap3__2487_ heichips25_sap3/net254 VPWR heichips25_sap3/_1900_ VGND heichips25_sap3/_1878_
+ heichips25_sap3/_1898_ sg13g2_o21ai_1
XFILLER_18_231 VPWR VGND sg13g2_decap_4
XFILLER_37_90 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3108_ heichips25_sap3/_0721_ heichips25_sap3/_0307_ heichips25_sap3/_0705_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__3039_ heichips25_sap3/net220 heichips25_sap3/_1778_ heichips25_sap3/_0649_
+ heichips25_sap3/_0652_ VPWR VGND sg13g2_nor3_1
Xheichips25_can_lehmann_fsm__2260_ heichips25_can_lehmann_fsm/net1181 VPWR heichips25_can_lehmann_fsm/_0578_
+ VGND heichips25_can_lehmann_fsm__2822_/Q heichips25_can_lehmann_fsm/_1044_ sg13g2_o21ai_1
XFILLER_30_996 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2191_ heichips25_can_lehmann_fsm/_1099_ heichips25_can_lehmann_fsm/net1192
+ heichips25_can_lehmann_fsm/_0524_ VPWR VGND sg13g2_nor2b_1
XFILLER_29_507 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1975_ heichips25_can_lehmann_fsm__2782_/Q heichips25_can_lehmann_fsm__2781_/Q
+ heichips25_can_lehmann_fsm/_1065_ heichips25_can_lehmann_fsm/_0334_ VPWR VGND sg13g2_nor3_1
XFILLER_17_27 VPWR VGND sg13g2_fill_2
Xheichips25_sap3_hold1224 heichips25_sap3__4043_/Q VPWR VGND heichips25_sap3/net1223
+ sg13g2_dlygate4sd3_1
XFILLER_33_790 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2527_ VGND VPWR heichips25_can_lehmann_fsm/_0916_ heichips25_can_lehmann_fsm/net415
+ heichips25_can_lehmann_fsm/_0163_ heichips25_can_lehmann_fsm/_0729_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2458_ heichips25_can_lehmann_fsm/net493 VPWR heichips25_can_lehmann_fsm/_0695_
+ VGND heichips25_can_lehmann_fsm__2904_/Q heichips25_can_lehmann_fsm/net405 sg13g2_o21ai_1
XFILLER_4_606 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2389_ VGND VPWR heichips25_can_lehmann_fsm/_0954_ heichips25_can_lehmann_fsm/net372
+ heichips25_can_lehmann_fsm/_0094_ heichips25_can_lehmann_fsm/_0660_ sg13g2_a21oi_1
Xclkbuf_4_0_0_heichips25_sap3\_sap_3_inst.alu_inst.clk clknet_0_heichips25_sap3\/sap_3_inst.alu_inst.clk
+ clknet_4_0_0_heichips25_sap3\/sap_3_inst.alu_inst.clk VPWR VGND sg13g2_buf_8
Xheichips25_sap3__2410_ heichips25_sap3/_1825_ heichips25_sap3/_1826_ heichips25_sap3/_1827_
+ VPWR VGND sg13g2_and2_1
Xheichips25_sap3__3390_ heichips25_sap3/_0965_ heichips25_sap3/_0991_ heichips25_sap3/_0998_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__2341_ heichips25_sap3/_1475_ heichips25_sap3/net225 heichips25_sap3/_1762_
+ VPWR VGND sg13g2_nor2_1
XFILLER_15_201 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2272_ heichips25_sap3/_1624_ heichips25_sap3/_1692_ heichips25_sap3/_1592_
+ heichips25_sap3/_1693_ VPWR VGND sg13g2_nand3_1
XFILLER_43_543 VPWR VGND sg13g2_fill_2
XFILLER_15_234 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__4011_ heichips25_sap3/net443 VGND VPWR heichips25_sap3/_0152_ heichips25_sap3__4011_/Q
+ clkload19/A sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2803__601 VPWR VGND net600 sg13g2_tiehi
XFILLER_30_248 VPWR VGND sg13g2_fill_2
XFILLER_7_499 VPWR VGND sg13g2_fill_2
XFILLER_7_488 VPWR VGND sg13g2_decap_8
XFILLER_48_1014 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__1987_ VPWR heichips25_sap3/_1413_ heichips25_sap3__4017_/Q VGND
+ sg13g2_inv_1
Xheichips25_sap3__3726_ heichips25_sap3__4026_/Q heichips25_sap3/net118 heichips25_sap3/_1244_
+ VPWR VGND sg13g2_nor2_1
XFILLER_2_182 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2853__790 VPWR VGND net789 sg13g2_tiehi
XFILLER_2_193 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3657_ heichips25_sap3/_1204_ heichips25_sap3/net119 uio_oe_sap3\[2\]
+ VPWR VGND sg13g2_nand2b_1
XFILLER_38_315 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3588_ heichips25_sap3/net120 VPWR heichips25_sap3/_1164_ VGND heichips25_sap3/net828
+ heichips25_sap3/_1144_ sg13g2_o21ai_1
Xheichips25_sap3__2608_ heichips25_sap3/_1635_ VPWR heichips25_sap3/_0279_ VGND heichips25_sap3/_1530_
+ heichips25_sap3/_1531_ sg13g2_o21ai_1
Xheichips25_sap3__2539_ heichips25_sap3/net286 heichips25_sap3/net289 heichips25_sap3/net279
+ heichips25_sap3/_0215_ VPWR VGND sg13g2_nor3_1
XFILLER_0_1027 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1760_ heichips25_can_lehmann_fsm/_1079_ heichips25_can_lehmann_fsm/_1032_
+ heichips25_can_lehmann_fsm__2799_/Q heichips25_can_lehmann_fsm/_1031_ heichips25_can_lehmann_fsm/net354
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2884__728 VPWR VGND net727 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__1691_ VPWR VGND heichips25_can_lehmann_fsm__3042_/Q heichips25_can_lehmann_fsm/_1014_
+ heichips25_can_lehmann_fsm/net331 heichips25_can_lehmann_fsm__2922_/Q heichips25_can_lehmann_fsm/_1015_
+ heichips25_can_lehmann_fsm/net313 sg13g2_a221oi_1
XFILLER_21_215 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2312_ heichips25_can_lehmann_fsm/_1052_ heichips25_can_lehmann_fsm/net206
+ heichips25_can_lehmann_fsm/_0620_ VPWR VGND heichips25_can_lehmann_fsm__2832_/Q
+ sg13g2_nand3b_1
Xheichips25_can_lehmann_fsm__2243_ VGND VPWR heichips25_can_lehmann_fsm/net205 heichips25_can_lehmann_fsm/_0563_
+ heichips25_can_lehmann_fsm/_0044_ heichips25_can_lehmann_fsm/_0564_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2174_ VGND VPWR heichips25_can_lehmann_fsm/_0508_ heichips25_can_lehmann_fsm/_0509_
+ heichips25_can_lehmann_fsm/_0029_ heichips25_can_lehmann_fsm/_0510_ sg13g2_a21oi_1
XFILLER_28_37 VPWR VGND sg13g2_fill_2
XFILLER_28_48 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1958_ heichips25_can_lehmann_fsm/net346 heichips25_can_lehmann_fsm/_1215_
+ heichips25_can_lehmann_fsm/_0320_ VPWR VGND sg13g2_nor2b_1
XFILLER_37_370 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2785__637 VPWR VGND net636 sg13g2_tiehi
Xheichips25_sap3_fanout443 heichips25_sap3/net446 heichips25_sap3/net443 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_hold1021 heichips25_sap3/_0017_ VPWR VGND heichips25_sap3/net1020
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__1889_ heichips25_can_lehmann_fsm/_1202_ heichips25_can_lehmann_fsm/net297
+ heichips25_can_lehmann_fsm__2911_/Q heichips25_can_lehmann_fsm/net314 heichips25_can_lehmann_fsm__2935_/Q
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3_fanout454 heichips25_sap3/net455 heichips25_sap3/net454 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_hold1032 heichips25_sap3__4039_/Q VPWR VGND heichips25_sap3/net1031
+ sg13g2_dlygate4sd3_1
XFILLER_40_557 VPWR VGND sg13g2_fill_2
Xheichips25_sap3_hold1065 heichips25_sap3__4058_/Q VPWR VGND heichips25_sap3/net1064
+ sg13g2_dlygate4sd3_1
XFILLER_21_771 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2890_ heichips25_sap3/_0504_ VPWR heichips25_sap3/_0531_ VGND heichips25_sap3/_0501_
+ heichips25_sap3/_0503_ sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm_fanout380 heichips25_can_lehmann_fsm/net388 heichips25_can_lehmann_fsm/net380
+ VPWR VGND sg13g2_buf_1
XFILLER_0_631 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3511_ VGND VPWR heichips25_sap3/_1380_ heichips25_sap3/net106 heichips25_sap3/_0090_
+ heichips25_sap3/_1105_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm_fanout391 heichips25_can_lehmann_fsm/net392 heichips25_can_lehmann_fsm/net391
+ VPWR VGND sg13g2_buf_1
Xheichips25_sap3__3442_ net47 heichips25_sap3/net68 heichips25_sap3/_1048_ VPWR VGND
+ sg13g2_nor2_1
Xheichips25_sap3__3373_ heichips25_sap3/net55 heichips25_sap3/_0980_ heichips25_sap3/_0981_
+ heichips25_sap3/_0982_ VPWR VGND sg13g2_nor3_1
Xheichips25_sap3__2324_ heichips25_sap3/_1694_ heichips25_sap3/_1712_ heichips25_sap3/_1731_
+ heichips25_sap3/_1745_ VPWR VGND sg13g2_nor3_1
Xheichips25_sap3__2255_ heichips25_sap3/_1661_ heichips25_sap3/_1673_ heichips25_sap3/_1675_
+ heichips25_sap3/_1676_ VPWR VGND sg13g2_nor3_1
Xheichips25_sap3__2186_ heichips25_sap3/_1468_ heichips25_sap3/_1547_ heichips25_sap3/_1607_
+ VPWR VGND sg13g2_nor2_1
XFILLER_16_587 VPWR VGND sg13g2_fill_2
XFILLER_34_80 VPWR VGND sg13g2_decap_8
XFILLER_11_281 VPWR VGND sg13g2_fill_1
XFILLER_7_285 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3709_ heichips25_sap3/_1114_ heichips25_sap3/_1237_ heichips25_sap3/_1238_
+ VPWR VGND sg13g2_and2_1
XFILLER_22_2 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2930_ net615 VGND VPWR heichips25_can_lehmann_fsm/_0155_
+ heichips25_can_lehmann_fsm__2930_/Q clknet_leaf_12_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2861_ net773 VGND VPWR heichips25_can_lehmann_fsm/net949
+ heichips25_can_lehmann_fsm__2861_/Q clknet_leaf_10_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1812_ heichips25_can_lehmann_fsm/_1128_ heichips25_can_lehmann_fsm/_1125_
+ heichips25_can_lehmann_fsm/_1126_ heichips25_can_lehmann_fsm/_1127_ VPWR VGND sg13g2_and3_1
Xheichips25_can_lehmann_fsm__2792_ net622 VGND VPWR heichips25_can_lehmann_fsm/net1228
+ heichips25_can_lehmann_fsm__2792_/Q clknet_leaf_1_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1743_ heichips25_can_lehmann_fsm/_1063_ heichips25_can_lehmann_fsm/_1062_
+ heichips25_can_lehmann_fsm__2779_/Q VPWR VGND sg13g2_nand2b_1
XFILLER_14_17 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1674_ heichips25_can_lehmann_fsm/net352 heichips25_can_lehmann_fsm/net353
+ heichips25_can_lehmann_fsm/_0998_ VPWR VGND sg13g2_nor2_1
Xheichips25_can_lehmann_fsm__2226_ heichips25_can_lehmann_fsm/_1105_ heichips25_can_lehmann_fsm/net1221
+ heichips25_can_lehmann_fsm/_0551_ VPWR VGND sg13g2_xor2_1
Xheichips25_can_lehmann_fsm__2157_ heichips25_can_lehmann_fsm/_0461_ heichips25_can_lehmann_fsm/_0493_
+ heichips25_can_lehmann_fsm/_0496_ VPWR VGND sg13g2_nor2_1
Xheichips25_can_lehmann_fsm__2088_ heichips25_can_lehmann_fsm__2799_/Q VPWR heichips25_can_lehmann_fsm/_0430_
+ VGND heichips25_can_lehmann_fsm/net345 heichips25_can_lehmann_fsm/_1056_ sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__3032__598 VPWR VGND net597 sg13g2_tiehi
XFILLER_18_819 VPWR VGND sg13g2_decap_4
XFILLER_29_167 VPWR VGND sg13g2_fill_2
XFILLER_26_841 VPWR VGND sg13g2_fill_1
XFILLER_44_159 VPWR VGND sg13g2_decap_4
XFILLER_44_148 VPWR VGND sg13g2_decap_4
Xheichips25_sap3_fanout240 heichips25_sap3/_1461_ heichips25_sap3/net240 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout273 heichips25_sap3__3923_/Q heichips25_sap3/net273 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3__2040_ heichips25_sap3/_1458_ heichips25_sap3/_1460_ heichips25_sap3/_1461_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3_fanout251 heichips25_sap3__4065_/Q heichips25_sap3/net251 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout262 heichips25_sap3/net263 heichips25_sap3/net262 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout284 heichips25_sap3/net285 heichips25_sap3/net284 VPWR VGND
+ sg13g2_buf_1
XFILLER_41_866 VPWR VGND sg13g2_fill_1
XFILLER_40_343 VPWR VGND sg13g2_decap_8
XFILLER_41_888 VPWR VGND sg13g2_fill_1
XFILLER_40_365 VPWR VGND sg13g2_decap_8
XFILLER_40_354 VPWR VGND sg13g2_fill_1
XFILLER_9_528 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3991_ heichips25_sap3/net459 VGND VPWR heichips25_sap3/_0132_ heichips25_sap3__3991_/Q
+ heichips25_sap3__3993_/CLK sg13g2_dfrbpq_1
Xheichips25_sap3__2942_ VGND VPWR heichips25_sap3/net65 heichips25_sap3/_0562_ heichips25_sap3/_0581_
+ heichips25_sap3/net203 sg13g2_a21oi_1
XFILLER_4_255 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2873_ heichips25_sap3/_0514_ VPWR heichips25_sap3/_0515_ VGND heichips25_sap3/net64
+ heichips25_sap3/_0513_ sg13g2_o21ai_1
XFILLER_45_1006 VPWR VGND sg13g2_fill_1
XFILLER_4_299 VPWR VGND sg13g2_decap_8
XFILLER_1_940 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__3015__763 VPWR VGND net762 sg13g2_tiehi
Xheichips25_sap3__3425_ heichips25_sap3/_1031_ heichips25_sap3/net104 heichips25_sap3__3946_/Q
+ heichips25_sap3/net110 heichips25_sap3__3954_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3356_ heichips25_sap3/_0965_ heichips25_sap3/_0959_ heichips25_sap3/_0964_
+ heichips25_sap3/net129 heichips25_sap3/_1400_ VPWR VGND sg13g2_a22oi_1
XFILLER_17_841 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2948__544 VPWR VGND net543 sg13g2_tiehi
Xheichips25_sap3__2307_ heichips25_sap3/_1599_ heichips25_sap3/net218 heichips25_sap3/_1726_
+ heichips25_sap3/_1727_ heichips25_sap3/_1728_ VPWR VGND sg13g2_nor4_1
Xheichips25_sap3__3287_ heichips25_sap3/_0777_ heichips25_sap3/net51 heichips25_sap3/_0899_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__2238_ heichips25_sap3/_1659_ heichips25_sap3/_1568_ heichips25_sap3/_1658_
+ VPWR VGND sg13g2_nand2_1
XFILLER_16_373 VPWR VGND sg13g2_fill_1
XFILLER_32_833 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2169_ heichips25_sap3/_1590_ heichips25_sap3/_1540_ heichips25_sap3/_1589_
+ VPWR VGND sg13g2_nand2_1
XFILLER_31_387 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__3060_ net653 VGND VPWR heichips25_can_lehmann_fsm/_0285_
+ heichips25_can_lehmann_fsm__3060_/Q clknet_leaf_14_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2011_ heichips25_can_lehmann_fsm__2779_/Q heichips25_can_lehmann_fsm/net191
+ heichips25_can_lehmann_fsm/_0365_ VPWR VGND sg13g2_nor2b_1
Xfanout507 net1 net507 VPWR VGND sg13g2_buf_1
XFILLER_6_1000 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2913_ net669 VGND VPWR heichips25_can_lehmann_fsm/_0138_
+ heichips25_can_lehmann_fsm__2913_/Q clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_39_465 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2844_ net807 VGND VPWR heichips25_can_lehmann_fsm/net852
+ heichips25_can_lehmann_fsm__2844_/Q clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_26_137 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2775_ net589 VGND VPWR heichips25_can_lehmann_fsm/_0000_
+ heichips25_can_lehmann_fsm__2775_/Q clknet_leaf_14_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2927__628 VPWR VGND net627 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__1726_ heichips25_can_lehmann_fsm/_1047_ heichips25_can_lehmann_fsm/_0973_
+ heichips25_can_lehmann_fsm/_1046_ VPWR VGND sg13g2_nand2_1
Xheichips25_can_lehmann_fsm__3027__667 VPWR VGND net666 sg13g2_tiehi
XFILLER_34_170 VPWR VGND sg13g2_fill_1
XFILLER_23_844 VPWR VGND sg13g2_fill_1
XFILLER_34_181 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__1657_ VPWR heichips25_can_lehmann_fsm/_0981_ heichips25_can_lehmann_fsm__2785_/Q
+ VGND sg13g2_inv_1
XFILLER_41_48 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1588_ VPWR heichips25_can_lehmann_fsm/_0912_ heichips25_can_lehmann_fsm/net904
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__2209_ heichips25_can_lehmann_fsm/_0538_ heichips25_can_lehmann_fsm/_1103_
+ heichips25_can_lehmann_fsm/_0537_ VPWR VGND sg13g2_nand2_1
XFILLER_2_737 VPWR VGND sg13g2_fill_2
XFILLER_1_214 VPWR VGND sg13g2_fill_1
XFILLER_1_269 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2910__676 VPWR VGND net675 sg13g2_tiehi
Xheichips25_sap3__3210_ heichips25_sap3/_0823_ heichips25_sap3/net138 heichips25_sap3__3979_/Q
+ heichips25_sap3/net140 heichips25_sap3__3987_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3141_ VPWR VGND heichips25_sap3/_0716_ heichips25_sap3/_0679_ heichips25_sap3/_0714_
+ heichips25_sap3/_0660_ heichips25_sap3/_0754_ heichips25_sap3/_0665_ sg13g2_a221oi_1
Xheichips25_sap3__3072_ heichips25_sap3/_1548_ VPWR heichips25_sap3/_0685_ VGND heichips25_sap3/_1464_
+ heichips25_sap3/_1552_ sg13g2_o21ai_1
XFILLER_14_800 VPWR VGND sg13g2_fill_2
XFILLER_26_671 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2023_ heichips25_sap3/net262 heichips25_sap3/net261 heichips25_sap3/_1444_
+ VPWR VGND heichips25_sap3/net264 sg13g2_nand3b_1
XFILLER_13_343 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_hold1160 heichips25_can_lehmann_fsm/_0056_ VPWR VGND heichips25_can_lehmann_fsm/net1159
+ sg13g2_dlygate4sd3_1
XFILLER_40_162 VPWR VGND sg13g2_fill_2
XFILLER_15_71 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm_hold1182 heichips25_can_lehmann_fsm__2823_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1181 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1193 heichips25_can_lehmann_fsm__2808_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1192 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1171 heichips25_can_lehmann_fsm__2827_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1170 sg13g2_dlygate4sd3_1
XFILLER_9_358 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3974_ heichips25_sap3/net457 VGND VPWR heichips25_sap3/_0115_ heichips25_sap3__3974_/Q
+ heichips25_sap3__3990_/CLK sg13g2_dfrbpq_1
Xheichips25_sap3__2925_ heichips25_sap3/_0338_ VPWR heichips25_sap3/_0564_ VGND heichips25_sap3/_0547_
+ heichips25_sap3/_0561_ sg13g2_o21ai_1
Xheichips25_sap3__2856_ heichips25_sap3/_0498_ heichips25_sap3/_0497_ heichips25_sap3/_0405_
+ VPWR VGND sg13g2_nand2b_1
Xheichips25_sap3_fanout90 heichips25_sap3/net92 heichips25_sap3/net90 VPWR VGND sg13g2_buf_1
Xheichips25_sap3__2787_ heichips25_sap3/_0432_ heichips25_sap3/_1452_ heichips25_sap3/_0431_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__3408_ VPWR heichips25_sap3/_1015_ heichips25_sap3/_1014_ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__2811__585 VPWR VGND net584 sg13g2_tiehi
XFILLER_36_457 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3339_ VPWR heichips25_sap3/_0949_ heichips25_sap3/_0948_ VGND sg13g2_inv_1
XFILLER_45_991 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2560_ heichips25_can_lehmann_fsm/net497 VPWR heichips25_can_lehmann_fsm/_0746_
+ VGND heichips25_can_lehmann_fsm__2954_/Q heichips25_can_lehmann_fsm/net386 sg13g2_o21ai_1
XFILLER_23_107 VPWR VGND sg13g2_fill_1
XFILLER_16_170 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2491_ VGND VPWR heichips25_can_lehmann_fsm/_0925_ heichips25_can_lehmann_fsm/net394
+ heichips25_can_lehmann_fsm/_0145_ heichips25_can_lehmann_fsm/_0711_ sg13g2_a21oi_1
XFILLER_20_847 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2996__626 VPWR VGND net625 sg13g2_tiehi
XFILLER_11_29 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__3043_ net710 VGND VPWR heichips25_can_lehmann_fsm/net878
+ heichips25_can_lehmann_fsm__3043_/Q clknet_leaf_21_clk sg13g2_dfrbpq_1
XFILLER_28_1012 VPWR VGND sg13g2_fill_2
XFILLER_39_284 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2827_ net552 VGND VPWR heichips25_can_lehmann_fsm/net1171
+ heichips25_can_lehmann_fsm__2827_/Q clknet_leaf_10_clk sg13g2_dfrbpq_1
XFILLER_14_107 VPWR VGND sg13g2_decap_8
XFILLER_14_129 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2758_ heichips25_can_lehmann_fsm/net488 VPWR heichips25_can_lehmann_fsm/_0845_
+ VGND heichips25_can_lehmann_fsm/net1084 heichips25_can_lehmann_fsm/net419 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2689_ VGND VPWR heichips25_can_lehmann_fsm/_0873_ heichips25_can_lehmann_fsm/net362
+ heichips25_can_lehmann_fsm/_0244_ heichips25_can_lehmann_fsm/_0810_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__1709_ VGND VPWR heichips25_can_lehmann_fsm/_1022_ heichips25_can_lehmann_fsm/_1028_
+ heichips25_can_lehmann_fsm/_1033_ heichips25_can_lehmann_fsm/_1032_ sg13g2_a21oi_1
XFILLER_6_317 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3690_ VGND VPWR heichips25_sap3/_1402_ heichips25_sap3/net113 heichips25_sap3/_0148_
+ heichips25_sap3/_1226_ sg13g2_a21oi_1
Xheichips25_sap3__2710_ VPWR heichips25_sap3/_0356_ heichips25_sap3/_0355_ VGND sg13g2_inv_1
Xheichips25_sap3__2641_ heichips25_sap3/_1544_ VPWR heichips25_sap3/_0308_ VGND heichips25_sap3/_0305_
+ heichips25_sap3/_0306_ sg13g2_o21ai_1
Xheichips25_sap3__2572_ heichips25_sap3/_0246_ heichips25_sap3__3891_/Q heichips25_sap3/_0243_
+ VPWR VGND sg13g2_nand2_1
XFILLER_46_755 VPWR VGND sg13g2_fill_1
XFILLER_45_298 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3124_ heichips25_sap3/_0732_ heichips25_sap3/net166 heichips25_sap3/_0737_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__3055_ VGND VPWR heichips25_sap3/_0668_ heichips25_sap3/_1725_ heichips25_sap3/_1363_
+ sg13g2_or2_1
Xheichips25_sap3__2006_ VPWR heichips25_sap3__4059_/D heichips25_sap3/net341 VGND
+ sg13g2_inv_1
XFILLER_13_173 VPWR VGND sg13g2_fill_2
XFILLER_13_184 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm_fanout209 heichips25_can_lehmann_fsm/net210 heichips25_can_lehmann_fsm/net209
+ VPWR VGND sg13g2_buf_1
Xheichips25_sap3__3957_ heichips25_sap3/net436 VGND VPWR heichips25_sap3/_0098_ heichips25_sap3__3957_/Q
+ heichips25_sap3__4005_/CLK sg13g2_dfrbpq_1
Xheichips25_sap3__2908_ heichips25_sap3/_0338_ heichips25_sap3/_0546_ heichips25_sap3/_0548_
+ VPWR VGND heichips25_sap3/_0547_ sg13g2_nand3b_1
XFILLER_5_394 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3888_ heichips25_sap3/net451 VGND VPWR heichips25_sap3/_0029_ heichips25_sap3__3888_/Q
+ heichips25_sap3__3921_/CLK sg13g2_dfrbpq_1
Xheichips25_sap3__2839_ heichips25_sap3/_0482_ heichips25_sap3/net285 heichips25_sap3/net212
+ VPWR VGND sg13g2_nand2_1
Xheichips25_can_lehmann_fsm__1991_ heichips25_can_lehmann_fsm/_0348_ heichips25_can_lehmann_fsm/net185
+ heichips25_can_lehmann_fsm/_0347_ heichips25_can_lehmann_fsm/net198 heichips25_can_lehmann_fsm__2783_/Q
+ VPWR VGND sg13g2_a22oi_1
XFILLER_37_711 VPWR VGND sg13g2_fill_2
XFILLER_36_276 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2612_ heichips25_can_lehmann_fsm/net485 VPWR heichips25_can_lehmann_fsm/_0772_
+ VGND heichips25_can_lehmann_fsm__2980_/Q heichips25_can_lehmann_fsm/net372 sg13g2_o21ai_1
Xclkbuf_leaf_16_clk clknet_2_2__leaf_clk clknet_leaf_16_clk VPWR VGND sg13g2_buf_8
Xheichips25_can_lehmann_fsm__2863__770 VPWR VGND net769 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2543_ VGND VPWR heichips25_can_lehmann_fsm/_0912_ heichips25_can_lehmann_fsm/net392
+ heichips25_can_lehmann_fsm/_0171_ heichips25_can_lehmann_fsm/_0737_ sg13g2_a21oi_1
XFILLER_32_460 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2474_ heichips25_can_lehmann_fsm/net483 VPWR heichips25_can_lehmann_fsm/_0703_
+ VGND heichips25_can_lehmann_fsm/net975 heichips25_can_lehmann_fsm/net415 sg13g2_o21ai_1
XFILLER_33_994 VPWR VGND sg13g2_fill_1
XFILLER_22_17 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2894__708 VPWR VGND net707 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__3026_ net674 VGND VPWR heichips25_can_lehmann_fsm/_0251_
+ heichips25_can_lehmann_fsm__3026_/Q clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_28_777 VPWR VGND sg13g2_fill_2
XFILLER_27_276 VPWR VGND sg13g2_decap_8
XFILLER_42_224 VPWR VGND sg13g2_fill_1
XFILLER_42_257 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm_hold843 heichips25_can_lehmann_fsm__3038_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net842 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold876 heichips25_can_lehmann_fsm/_0190_ VPWR VGND heichips25_can_lehmann_fsm/net875
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold854 heichips25_can_lehmann_fsm__3015_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net853 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold865 heichips25_can_lehmann_fsm/_0159_ VPWR VGND heichips25_can_lehmann_fsm/net864
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold887 heichips25_can_lehmann_fsm/_0192_ VPWR VGND heichips25_can_lehmann_fsm/net886
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold898 heichips25_can_lehmann_fsm__2978_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net897 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__2795__617 VPWR VGND net616 sg13g2_tiehi
Xheichips25_sap3__3811_ heichips25_sap3/net340 heichips25_sap3/net891 heichips25_sap3/_1318_
+ heichips25_sap3/_0177_ VPWR VGND sg13g2_a21o_1
XFILLER_10_198 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3742_ VGND VPWR heichips25_sap3/_0289_ heichips25_sap3/_1246_ heichips25_sap3/_0171_
+ heichips25_sap3/net1163 sg13g2_a21oi_1
XFILLER_3_854 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3673_ heichips25_sap3/_1216_ heichips25_sap3/_0992_ heichips25_sap3/_1015_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__2624_ heichips25_sap3/_0292_ heichips25_sap3/_1682_ heichips25_sap3/_1537_
+ heichips25_sap3/_1627_ heichips25_sap3/_1513_ VPWR VGND sg13g2_a22oi_1
X_10_ uo_out_fsm\[4\] uo_out_sap3\[4\] net507 net39 VPWR VGND sg13g2_mux2_1
Xheichips25_sap3__2555_ heichips25_sap3/_0230_ heichips25_sap3/net71 heichips25_sap3__3974_/Q
+ heichips25_sap3/net87 heichips25_sap3__3942_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_19_8 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2486_ heichips25_sap3/_1878_ heichips25_sap3/_1898_ heichips25_sap3/_1899_
+ VPWR VGND sg13g2_nor2_1
XFILLER_34_714 VPWR VGND sg13g2_decap_8
XFILLER_34_736 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3107_ heichips25_sap3/_0720_ heichips25_sap3/_0680_ heichips25_sap3/net152
+ VPWR VGND sg13g2_nand2_1
XFILLER_14_471 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3038_ VPWR VGND heichips25_sap3/_1664_ heichips25_sap3/_0648_ heichips25_sap3/_0650_
+ heichips25_sap3/net263 heichips25_sap3/_0651_ heichips25_sap3/_1773_ sg13g2_a221oi_1
Xheichips25_can_lehmann_fsm__2190_ VGND VPWR heichips25_can_lehmann_fsm/net160 heichips25_can_lehmann_fsm/_0522_
+ heichips25_can_lehmann_fsm/_0032_ heichips25_can_lehmann_fsm/_0523_ sg13g2_a21oi_1
Xclkbuf_leaf_5_clk clknet_2_1__leaf_clk clknet_leaf_5_clk VPWR VGND sg13g2_buf_8
XFILLER_38_0 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__3030__630 VPWR VGND net629 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__1974_ VGND VPWR heichips25_can_lehmann_fsm/net1248 heichips25_can_lehmann_fsm/net190
+ heichips25_can_lehmann_fsm/_0333_ heichips25_can_lehmann_fsm/net196 sg13g2_a21oi_1
XFILLER_37_541 VPWR VGND sg13g2_decap_8
Xheichips25_sap3_hold1225 heichips25_sap3__4042_/Q VPWR VGND heichips25_sap3/net1224
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__2526_ heichips25_can_lehmann_fsm/net483 VPWR heichips25_can_lehmann_fsm/_0729_
+ VGND heichips25_can_lehmann_fsm__2938_/Q heichips25_can_lehmann_fsm/net415 sg13g2_o21ai_1
XFILLER_33_780 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2457_ VGND VPWR heichips25_can_lehmann_fsm/_0933_ heichips25_can_lehmann_fsm/net365
+ heichips25_can_lehmann_fsm/_0128_ heichips25_can_lehmann_fsm/_0694_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2388_ heichips25_can_lehmann_fsm/net480 VPWR heichips25_can_lehmann_fsm/_0660_
+ VGND heichips25_can_lehmann_fsm__2868_/Q heichips25_can_lehmann_fsm/net372 sg13g2_o21ai_1
XFILLER_0_824 VPWR VGND sg13g2_fill_2
XFILLER_0_846 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__3009_ net810 VGND VPWR heichips25_can_lehmann_fsm/net868
+ heichips25_can_lehmann_fsm__3009_/Q clknet_leaf_17_clk sg13g2_dfrbpq_1
Xclkbuf_5_16__f_heichips25_sap3\_sap_3_inst.alu_inst.clk clkload23/A clknet_4_8_0_heichips25_sap3\/sap_3_inst.alu_inst.clk
+ VPWR VGND sg13g2_buf_16
Xheichips25_sap3__2340_ heichips25_sap3/_1515_ heichips25_sap3/_1605_ heichips25_sap3/net264
+ heichips25_sap3/_1761_ VPWR VGND sg13g2_nand3_1
Xheichips25_sap3__2271_ heichips25_sap3/_1540_ VPWR heichips25_sap3/_1692_ VGND heichips25_sap3/_1538_
+ heichips25_sap3/_1691_ sg13g2_o21ai_1
Xheichips25_sap3__4010_ heichips25_sap3/net445 VGND VPWR heichips25_sap3/_0151_ heichips25_sap3__4010_/Q
+ clkload22/A sg13g2_dfrbpq_1
XFILLER_43_533 VPWR VGND sg13g2_fill_2
XFILLER_15_213 VPWR VGND sg13g2_decap_4
XFILLER_43_566 VPWR VGND sg13g2_decap_8
XFILLER_12_953 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__1986_ VPWR heichips25_sap3/_1412_ heichips25_sap3__3937_/Q VGND
+ sg13g2_inv_1
Xheichips25_sap3__3725_ heichips25_sap3__4025_/Q heichips25_sap3/_1141_ heichips25_sap3/net118
+ heichips25_sap3/_0166_ VPWR VGND sg13g2_mux2_1
XFILLER_3_662 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3656_ heichips25_sap3/_0889_ heichips25_sap3/_1202_ heichips25_sap3/_1203_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__2607_ heichips25_sap3/_0278_ heichips25_sap3/_1636_ heichips25_sap3/_1553_
+ VPWR VGND sg13g2_nand2b_1
Xheichips25_sap3__3587_ heichips25_sap3/_1160_ heichips25_sap3/_1163_ heichips25_sap3/_0108_
+ VPWR VGND sg13g2_nor2b_1
Xheichips25_sap3__2538_ heichips25_sap3/_1886_ heichips25_sap3/_0213_ heichips25_sap3/_0214_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__2469_ heichips25_sap3/_1882_ heichips25_sap3/_1434_ heichips25_sap3/_1782_
+ VPWR VGND sg13g2_nand2_1
XFILLER_0_1006 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1690_ heichips25_can_lehmann_fsm/_1012_ heichips25_can_lehmann_fsm/_1013_
+ heichips25_can_lehmann_fsm/_1011_ heichips25_can_lehmann_fsm/_1014_ VPWR VGND sg13g2_nand3_1
XFILLER_9_51 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2311_ VGND VPWR heichips25_can_lehmann_fsm/net206 heichips25_can_lehmann_fsm/net1189
+ heichips25_can_lehmann_fsm/_0057_ heichips25_can_lehmann_fsm/_0619_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2242_ heichips25_can_lehmann_fsm/net329 VPWR heichips25_can_lehmann_fsm/_0564_
+ VGND heichips25_can_lehmann_fsm/net1174 heichips25_can_lehmann_fsm/net205 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2173_ heichips25_can_lehmann_fsm/net325 VPWR heichips25_can_lehmann_fsm/_0510_
+ VGND heichips25_can_lehmann_fsm/net1215 heichips25_can_lehmann_fsm/net160 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__1957_ heichips25_can_lehmann_fsm/net321 VPWR heichips25_can_lehmann_fsm/_0319_
+ VGND heichips25_can_lehmann_fsm/net1253 heichips25_can_lehmann_fsm/net178 sg13g2_o21ai_1
Xheichips25_sap3_fanout433 heichips25_sap3/net437 heichips25_sap3/net433 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout444 heichips25_sap3/net445 heichips25_sap3/net444 VPWR VGND
+ sg13g2_buf_1
Xheichips25_can_lehmann_fsm__1888_ heichips25_can_lehmann_fsm/_1201_ heichips25_can_lehmann_fsm/net307
+ heichips25_can_lehmann_fsm__2959_/Q heichips25_can_lehmann_fsm/net311 heichips25_can_lehmann_fsm__3031_/Q
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3_fanout455 heichips25_sap3/net463 heichips25_sap3/net455 VPWR VGND
+ sg13g2_buf_1
XFILLER_25_566 VPWR VGND sg13g2_decap_4
Xheichips25_sap3_hold1033 heichips25_sap3/_0180_ VPWR VGND heichips25_sap3/net1032
+ sg13g2_dlygate4sd3_1
XFILLER_12_216 VPWR VGND sg13g2_decap_8
Xheichips25_sap3_hold1066 heichips25_sap3/_0287_ VPWR VGND heichips25_sap3/net1065
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__2941__572 VPWR VGND net571 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2509_ VGND VPWR heichips25_can_lehmann_fsm/_0920_ heichips25_can_lehmann_fsm/net381
+ heichips25_can_lehmann_fsm/_0154_ heichips25_can_lehmann_fsm/_0720_ sg13g2_a21oi_1
XFILLER_5_938 VPWR VGND sg13g2_fill_2
XFILLER_4_459 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm_fanout370 heichips25_can_lehmann_fsm/net371 heichips25_can_lehmann_fsm/net370
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout392 heichips25_can_lehmann_fsm/net393 heichips25_can_lehmann_fsm/net392
+ VPWR VGND sg13g2_buf_1
Xheichips25_sap3__3510_ VPWR VGND heichips25_sap3/_1103_ heichips25_sap3/net106 heichips25_sap3/_1100_
+ heichips25_sap3/net97 heichips25_sap3/_1105_ heichips25_sap3/_0928_ sg13g2_a221oi_1
Xheichips25_can_lehmann_fsm_fanout381 heichips25_can_lehmann_fsm/net388 heichips25_can_lehmann_fsm/net381
+ VPWR VGND sg13g2_buf_1
Xheichips25_sap3__3441_ VPWR heichips25_sap3/_1047_ heichips25_sap3/_1046_ VGND sg13g2_inv_1
Xheichips25_sap3__3372_ net46 uio_oe_sap3\[4\] heichips25_sap3/net68 heichips25_sap3/_0981_
+ VPWR VGND sg13g2_mux2_1
Xheichips25_sap3__2323_ heichips25_sap3/_1680_ heichips25_sap3/_1736_ heichips25_sap3/_1744_
+ VPWR VGND sg13g2_and2_1
XFILLER_16_511 VPWR VGND sg13g2_decap_4
XFILLER_28_382 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2254_ heichips25_sap3/_1667_ heichips25_sap3/_1674_ heichips25_sap3/_1665_
+ heichips25_sap3/_1675_ VPWR VGND sg13g2_nand3_1
Xheichips25_sap3__2185_ heichips25_sap3/_1606_ heichips25_sap3/_1459_ heichips25_sap3/_1477_
+ VPWR VGND sg13g2_nand2_1
XFILLER_31_525 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2920__656 VPWR VGND net655 sg13g2_tiehi
Xheichips25_sap3__3708_ uio_oe_sap3\[4\] heichips25_sap3/net114 heichips25_sap3/_1237_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__1969_ VPWR heichips25_sap3/_1395_ heichips25_sap3__3955_/Q VGND
+ sg13g2_inv_1
XFILLER_3_492 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3639_ heichips25_sap3/_1138_ heichips25_sap3__3991_/Q heichips25_sap3/net93
+ heichips25_sap3/_0132_ VPWR VGND sg13g2_mux2_1
XFILLER_38_102 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2860_ net775 VGND VPWR heichips25_can_lehmann_fsm/_0085_
+ heichips25_can_lehmann_fsm__2860_/Q clknet_leaf_10_clk sg13g2_dfrbpq_1
XFILLER_38_179 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1811_ heichips25_can_lehmann_fsm/_1127_ heichips25_can_lehmann_fsm/net305
+ heichips25_can_lehmann_fsm__2947_/Q heichips25_can_lehmann_fsm/net310 heichips25_can_lehmann_fsm__3019_/Q
+ VPWR VGND sg13g2_a22oi_1
XFILLER_26_308 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2791_ net624 VGND VPWR heichips25_can_lehmann_fsm/net1239
+ heichips25_can_lehmann_fsm__2791_/Q clknet_leaf_1_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1742_ heichips25_can_lehmann_fsm__2778_/Q heichips25_can_lehmann_fsm/_1061_
+ heichips25_can_lehmann_fsm/_1062_ VPWR VGND sg13g2_nor2b_1
XFILLER_19_360 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1673_ heichips25_can_lehmann_fsm/net348 heichips25_can_lehmann_fsm/_0996_
+ heichips25_can_lehmann_fsm/_0997_ VPWR VGND sg13g2_nor2_1
Xheichips25_can_lehmann_fsm__2999__602 VPWR VGND net601 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2821__565 VPWR VGND net564 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2225_ VGND VPWR heichips25_can_lehmann_fsm/net161 heichips25_can_lehmann_fsm/_0549_
+ heichips25_can_lehmann_fsm/_0040_ heichips25_can_lehmann_fsm/_0550_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2156_ heichips25_can_lehmann_fsm/_0492_ heichips25_can_lehmann_fsm/net205
+ heichips25_can_lehmann_fsm/_0461_ heichips25_can_lehmann_fsm/_0495_ VPWR VGND sg13g2_a21o_1
Xheichips25_can_lehmann_fsm__2087_ VGND VPWR heichips25_can_lehmann_fsm/_0426_ heichips25_can_lehmann_fsm/_0428_
+ heichips25_can_lehmann_fsm/_0023_ heichips25_can_lehmann_fsm/_0429_ sg13g2_a21oi_1
XFILLER_44_138 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2989_ net668 VGND VPWR heichips25_can_lehmann_fsm/_0214_
+ heichips25_can_lehmann_fsm__2989_/Q clknet_leaf_18_clk sg13g2_dfrbpq_1
Xheichips25_sap3_fanout230 heichips25_sap3/_1479_ heichips25_sap3/net230 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout241 heichips25_sap3/_1452_ heichips25_sap3/net241 VPWR VGND
+ sg13g2_buf_1
XFILLER_40_300 VPWR VGND sg13g2_decap_8
Xheichips25_sap3_fanout263 heichips25_sap3__3927_/Q heichips25_sap3/net263 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout252 heichips25_sap3__4064_/Q heichips25_sap3/net252 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout274 heichips25_sap3__3906_/Q heichips25_sap3/net274 VPWR VGND
+ sg13g2_buf_1
XFILLER_26_897 VPWR VGND sg13g2_fill_2
XFILLER_40_322 VPWR VGND sg13g2_fill_2
Xheichips25_sap3_fanout285 heichips25_sap3__3901_/Q heichips25_sap3/net285 VPWR VGND
+ sg13g2_buf_1
XFILLER_41_878 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3990_ heichips25_sap3/net457 VGND VPWR heichips25_sap3/_0131_ heichips25_sap3__3990_/Q
+ heichips25_sap3__3990_/CLK sg13g2_dfrbpq_1
Xheichips25_sap3__2941_ heichips25_sap3/_0574_ VPWR heichips25_sap3/_0580_ VGND heichips25_sap3/_1869_
+ heichips25_sap3/_0579_ sg13g2_o21ai_1
Xheichips25_sap3__2872_ VGND VPWR heichips25_sap3/_0378_ heichips25_sap3/net64 heichips25_sap3/_0514_
+ heichips25_sap3/net203 sg13g2_a21oi_1
XFILLER_4_234 VPWR VGND sg13g2_fill_1
XFILLER_49_901 VPWR VGND sg13g2_fill_2
XFILLER_0_473 VPWR VGND sg13g2_decap_8
XFILLER_1_996 VPWR VGND sg13g2_decap_8
XFILLER_49_967 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3424_ VPWR VGND heichips25_sap3__4002_/Q heichips25_sap3/net124
+ heichips25_sap3/net146 heichips25_sap3__4018_/Q heichips25_sap3/_1030_ heichips25_sap3/net118
+ sg13g2_a221oi_1
XFILLER_0_484 VPWR VGND sg13g2_fill_2
XFILLER_49_989 VPWR VGND sg13g2_decap_8
XFILLER_36_606 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3355_ VPWR VGND heichips25_sap3__3943_/Q heichips25_sap3/_0963_
+ heichips25_sap3/net104 heichips25_sap3__3951_/Q heichips25_sap3/_0964_ heichips25_sap3/net109
+ sg13g2_a221oi_1
Xheichips25_sap3__2306_ heichips25_sap3/_1462_ heichips25_sap3/_1518_ heichips25_sap3/_1727_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__3286_ heichips25_sap3/_0898_ heichips25_sap3/_0895_ heichips25_sap3/_0897_
+ heichips25_sap3/net128 heichips25_sap3/_1385_ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2237_ heichips25_sap3/_1527_ heichips25_sap3/_1565_ heichips25_sap3/_1504_
+ heichips25_sap3/_1658_ VPWR VGND sg13g2_nand3_1
XFILLER_16_363 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2168_ heichips25_sap3/_1564_ heichips25_sap3/_1588_ heichips25_sap3/_1556_
+ heichips25_sap3/_1589_ VPWR VGND sg13g2_nand3_1
XFILLER_31_355 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2099_ heichips25_sap3/net256 heichips25_sap3/_1446_ heichips25_sap3/_1506_
+ heichips25_sap3/_1520_ VPWR VGND sg13g2_nor3_1
XFILLER_6_41 VPWR VGND sg13g2_decap_8
XFILLER_8_595 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2010_ heichips25_can_lehmann_fsm/_0364_ heichips25_can_lehmann_fsm/net184
+ heichips25_can_lehmann_fsm/_0363_ VPWR VGND sg13g2_nand2_1
XFILLER_6_1012 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2912_ net671 VGND VPWR heichips25_can_lehmann_fsm/_0137_
+ heichips25_can_lehmann_fsm__2912_/Q clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_27_617 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2843_ net809 VGND VPWR heichips25_can_lehmann_fsm/_0068_
+ heichips25_can_lehmann_fsm__2843_/Q clknet_leaf_4_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2774_ VGND VPWR heichips25_can_lehmann_fsm/_1041_ heichips25_can_lehmann_fsm/_1042_
+ heichips25_can_lehmann_fsm/_0288_ heichips25_can_lehmann_fsm/_1176_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__1725_ heichips25_can_lehmann_fsm__2824_/Q heichips25_can_lehmann_fsm__2823_/Q
+ heichips25_can_lehmann_fsm__2822_/Q heichips25_can_lehmann_fsm/_1044_ heichips25_can_lehmann_fsm/_1046_
+ VPWR VGND sg13g2_nor4_1
XFILLER_22_300 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1656_ VPWR heichips25_can_lehmann_fsm/_0980_ heichips25_can_lehmann_fsm__2790_/Q
+ VGND sg13g2_inv_1
XFILLER_22_355 VPWR VGND sg13g2_decap_8
XFILLER_22_366 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1587_ VPWR heichips25_can_lehmann_fsm/_0911_ heichips25_can_lehmann_fsm/net934
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__2208_ heichips25_can_lehmann_fsm/net1207 VPWR heichips25_can_lehmann_fsm/_0537_
+ VGND heichips25_can_lehmann_fsm__2811_/Q heichips25_can_lehmann_fsm/_1102_ sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2873__750 VPWR VGND net749 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2139_ heichips25_can_lehmann_fsm/_0478_ heichips25_can_lehmann_fsm/net308
+ heichips25_can_lehmann_fsm__2956_/Q heichips25_can_lehmann_fsm/net319 heichips25_can_lehmann_fsm__3004_/Q
+ VPWR VGND sg13g2_a22oi_1
XFILLER_17_116 VPWR VGND sg13g2_decap_8
XFILLER_17_127 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3140_ heichips25_sap3/_0753_ heichips25_sap3/_0717_ heichips25_sap3/net150
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__3071_ heichips25_sap3/net228 heichips25_sap3/_1668_ heichips25_sap3/_1474_
+ heichips25_sap3/_0684_ VPWR VGND sg13g2_nand3_1
Xheichips25_sap3__2022_ heichips25_sap3/net265 heichips25_sap3/net256 heichips25_sap3/_1443_
+ VPWR VGND sg13g2_nor2_1
XFILLER_13_311 VPWR VGND sg13g2_decap_8
XFILLER_26_694 VPWR VGND sg13g2_fill_1
XFILLER_9_315 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm_hold1183 heichips25_can_lehmann_fsm__2825_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1182 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1172 heichips25_can_lehmann_fsm/_0052_ VPWR VGND heichips25_can_lehmann_fsm/net1171
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1161 heichips25_can_lehmann_fsm__3034_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1160 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1194 heichips25_can_lehmann_fsm/_0033_ VPWR VGND heichips25_can_lehmann_fsm/net1193
+ sg13g2_dlygate4sd3_1
Xheichips25_sap3__3973_ heichips25_sap3/net447 VGND VPWR heichips25_sap3/_0114_ heichips25_sap3__3973_/Q
+ heichips25_sap3__4003_/CLK sg13g2_dfrbpq_1
Xheichips25_sap3_hold892 heichips25_sap3__4036_/Q VPWR VGND heichips25_sap3/net891
+ sg13g2_dlygate4sd3_1
Xheichips25_sap3__2924_ heichips25_sap3/_0563_ heichips25_sap3/_0547_ heichips25_sap3/_0561_
+ VPWR VGND sg13g2_nand2_1
XFILLER_12_1028 VPWR VGND sg13g2_fill_1
XFILLER_5_554 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2855_ heichips25_sap3/_0404_ VPWR heichips25_sap3/_0497_ VGND heichips25_sap3/_0402_
+ heichips25_sap3/_0403_ sg13g2_o21ai_1
Xheichips25_sap3_fanout80 heichips25_sap3/_1741_ heichips25_sap3/net80 VPWR VGND sg13g2_buf_1
Xheichips25_sap3_fanout91 heichips25_sap3/net92 heichips25_sap3/net91 VPWR VGND sg13g2_buf_1
Xheichips25_sap3__2786_ heichips25_sap3/_1767_ heichips25_sap3/_0430_ heichips25_sap3/net221
+ heichips25_sap3/_0431_ VPWR VGND sg13g2_nand3_1
XFILLER_49_786 VPWR VGND sg13g2_decap_8
XFILLER_48_263 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3407_ heichips25_sap3/_1014_ heichips25_sap3/_1008_ heichips25_sap3/_1013_
+ heichips25_sap3/net126 heichips25_sap3/_1412_ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3338_ heichips25_sap3/net98 VPWR heichips25_sap3/_0948_ VGND heichips25_sap3/net128
+ heichips25_sap3/_0947_ sg13g2_o21ai_1
Xheichips25_sap3__3269_ VPWR heichips25_sap3/_0882_ heichips25_sap3/net131 VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__2490_ heichips25_can_lehmann_fsm/net464 VPWR heichips25_can_lehmann_fsm/_0711_
+ VGND heichips25_can_lehmann_fsm__2920_/Q heichips25_can_lehmann_fsm/net394 sg13g2_o21ai_1
XFILLER_31_152 VPWR VGND sg13g2_decap_8
XFILLER_31_163 VPWR VGND sg13g2_fill_1
XFILLER_9_871 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__3042_ net726 VGND VPWR heichips25_can_lehmann_fsm/_0267_
+ heichips25_can_lehmann_fsm__3042_/Q clknet_leaf_21_clk sg13g2_dfrbpq_1
XFILLER_28_1024 VPWR VGND sg13g2_decap_4
XFILLER_39_274 VPWR VGND sg13g2_decap_4
XFILLER_27_403 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2826_ net554 VGND VPWR heichips25_can_lehmann_fsm/_0051_
+ heichips25_can_lehmann_fsm__2826_/Q clknet_leaf_10_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2757_ VGND VPWR heichips25_can_lehmann_fsm/_0855_ heichips25_can_lehmann_fsm/net384
+ heichips25_can_lehmann_fsm/_0278_ heichips25_can_lehmann_fsm/_0844_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2688_ heichips25_can_lehmann_fsm/net468 VPWR heichips25_can_lehmann_fsm/_0810_
+ VGND heichips25_can_lehmann_fsm__3018_/Q heichips25_can_lehmann_fsm/net359 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__1708_ heichips25_can_lehmann_fsm/_1010_ heichips25_can_lehmann_fsm/_1030_
+ heichips25_can_lehmann_fsm/_1032_ VPWR VGND sg13g2_and2_1
Xheichips25_can_lehmann_fsm__1639_ VPWR heichips25_can_lehmann_fsm/_0963_ heichips25_can_lehmann_fsm/net840
+ VGND sg13g2_inv_1
Xheichips25_sap3__2640_ VGND VPWR heichips25_sap3/net236 heichips25_sap3/_1543_ heichips25_sap3/_0307_
+ heichips25_sap3/_1532_ sg13g2_a21oi_1
Xheichips25_sap3__2571_ heichips25_sap3/_0244_ VPWR heichips25_sap3/_0245_ VGND heichips25_sap3/net275
+ heichips25_sap3/_1801_ sg13g2_o21ai_1
XFILLER_18_403 VPWR VGND sg13g2_fill_1
XFILLER_19_948 VPWR VGND sg13g2_fill_2
XFILLER_34_929 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3123_ heichips25_sap3/_0734_ heichips25_sap3/_0735_ heichips25_sap3/_0733_
+ heichips25_sap3/_0736_ VPWR VGND sg13g2_nand3_1
XFILLER_26_82 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3054_ heichips25_sap3/_0659_ heichips25_sap3/net241 heichips25_sap3/_0664_
+ heichips25_sap3/_0667_ VPWR VGND sg13g2_a21o_1
XFILLER_9_101 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2005_ VPWR heichips25_sap3/_1430_ heichips25_sap3__4072_/A VGND
+ sg13g2_inv_1
XFILLER_9_189 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3956_ heichips25_sap3/net434 VGND VPWR heichips25_sap3/_0097_ heichips25_sap3__3956_/Q
+ heichips25_sap3__4012_/CLK sg13g2_dfrbpq_1
Xheichips25_sap3__3887_ heichips25_sap3/net451 VGND VPWR heichips25_sap3/_0028_ heichips25_sap3__3887_/Q
+ heichips25_sap3__3921_/CLK sg13g2_dfrbpq_1
XFILLER_5_351 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2907_ heichips25_sap3/_0379_ heichips25_sap3/_0522_ heichips25_sap3/_0545_
+ heichips25_sap3/_0547_ VPWR VGND sg13g2_nor3_1
Xheichips25_sap3__2838_ heichips25_sap3/_0481_ heichips25_sap3/_0417_ heichips25_sap3/net287
+ heichips25_sap3/_0416_ heichips25_sap3/net282 VPWR VGND sg13g2_a22oi_1
XFILLER_3_42 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2769_ VGND VPWR heichips25_sap3/net274 heichips25_sap3/_1399_ heichips25_sap3/_0415_
+ heichips25_sap3/_0414_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__1990_ heichips25_can_lehmann_fsm/_1067_ VPWR heichips25_can_lehmann_fsm/_0347_
+ VGND heichips25_can_lehmann_fsm/_0982_ heichips25_can_lehmann_fsm/_0339_ sg13g2_o21ai_1
XFILLER_3_1026 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2611_ VGND VPWR heichips25_can_lehmann_fsm/_0895_ heichips25_can_lehmann_fsm/net425
+ heichips25_can_lehmann_fsm/_0205_ heichips25_can_lehmann_fsm/_0771_ sg13g2_a21oi_1
XFILLER_36_299 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__3063__687 VPWR VGND net686 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2542_ heichips25_can_lehmann_fsm/net467 VPWR heichips25_can_lehmann_fsm/_0737_
+ VGND heichips25_can_lehmann_fsm__2946_/Q heichips25_can_lehmann_fsm/net392 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2473_ VGND VPWR heichips25_can_lehmann_fsm/_0929_ heichips25_can_lehmann_fsm/net376
+ heichips25_can_lehmann_fsm/_0136_ heichips25_can_lehmann_fsm/_0702_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__3025_ net682 VGND VPWR heichips25_can_lehmann_fsm/net1075
+ heichips25_can_lehmann_fsm__3025_/Q clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_27_233 VPWR VGND sg13g2_fill_2
XFILLER_42_203 VPWR VGND sg13g2_decap_8
XFILLER_27_255 VPWR VGND sg13g2_decap_8
XFILLER_28_789 VPWR VGND sg13g2_fill_2
XFILLER_43_737 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2809_ net588 VGND VPWR heichips25_can_lehmann_fsm/net1199
+ heichips25_can_lehmann_fsm__2809_/Q clknet_leaf_5_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__3042__727 VPWR VGND net726 sg13g2_tiehi
XFILLER_24_962 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm_hold844 heichips25_can_lehmann_fsm/_0264_ VPWR VGND heichips25_can_lehmann_fsm/net843
+ sg13g2_dlygate4sd3_1
XFILLER_10_100 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm_hold877 heichips25_can_lehmann_fsm__2896_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net876 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold866 heichips25_can_lehmann_fsm__2895_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net865 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold855 heichips25_can_lehmann_fsm/_0241_ VPWR VGND heichips25_can_lehmann_fsm/net854
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold899 heichips25_can_lehmann_fsm__2853_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net898 sg13g2_dlygate4sd3_1
XFILLER_6_104 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm_hold888 heichips25_can_lehmann_fsm__2969_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net887 sg13g2_dlygate4sd3_1
Xheichips25_sap3__3810_ VPWR VGND heichips25_sap3/_1317_ heichips25_sap3/net340 heichips25_sap3/_1311_
+ heichips25_sap3/_1400_ heichips25_sap3/_1318_ heichips25_sap3/net291 sg13g2_a221oi_1
XFILLER_12_51 VPWR VGND sg13g2_fill_2
XFILLER_12_62 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3741_ VGND VPWR heichips25_sap3__4029_/Q heichips25_sap3/_1246_
+ heichips25_sap3/_1255_ heichips25_sap3/net1162 sg13g2_a21oi_1
XFILLER_3_800 VPWR VGND sg13g2_fill_1
XFILLER_12_95 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3672_ heichips25_sap3/_0141_ heichips25_sap3/_1121_ heichips25_sap3/_1215_
+ heichips25_sap3/net111 heichips25_sap3/_1407_ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2623_ heichips25_sap3/_0000_ heichips25_sap3/net1131 heichips25_sap3/net832
+ VPWR VGND sg13g2_nand2b_1
Xheichips25_sap3__2554_ heichips25_sap3/_0229_ heichips25_sap3/net76 heichips25_sap3__3982_/Q
+ heichips25_sap3/net216 heichips25_sap3__4006_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2485_ heichips25_sap3/_1885_ heichips25_sap3/_1887_ heichips25_sap3/_1888_
+ heichips25_sap3/_1897_ heichips25_sap3/_1898_ VPWR VGND sg13g2_and4_1
XFILLER_18_211 VPWR VGND sg13g2_decap_8
XFILLER_19_756 VPWR VGND sg13g2_fill_2
XFILLER_19_767 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__3047__638 VPWR VGND net637 sg13g2_tiehi
XFILLER_18_299 VPWR VGND sg13g2_decap_8
XFILLER_14_450 VPWR VGND sg13g2_decap_8
XFILLER_15_951 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3106_ heichips25_sap3/_0680_ heichips25_sap3/net152 heichips25_sap3/_0719_
+ VPWR VGND sg13g2_and2_1
XFILLER_33_247 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3037_ heichips25_sap3/_0650_ heichips25_sap3/_1486_ heichips25_sap3/_1625_
+ VPWR VGND sg13g2_nand2_1
XFILLER_30_976 VPWR VGND sg13g2_decap_8
XFILLER_6_693 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3939_ heichips25_sap3/net456 VGND VPWR heichips25_sap3/_0080_ heichips25_sap3__3939_/Q
+ clkload28/A sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1973_ VGND VPWR heichips25_can_lehmann_fsm/_0330_ heichips25_can_lehmann_fsm/_0331_
+ heichips25_can_lehmann_fsm/_0006_ heichips25_can_lehmann_fsm/_0332_ sg13g2_a21oi_1
XFILLER_37_564 VPWR VGND sg13g2_decap_8
Xheichips25_sap3_hold1226 heichips25_sap3__4058_/Q VPWR VGND heichips25_sap3/net1225
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__2525_ VGND VPWR heichips25_can_lehmann_fsm/_0916_ heichips25_can_lehmann_fsm/net375
+ heichips25_can_lehmann_fsm/_0162_ heichips25_can_lehmann_fsm/_0728_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2456_ heichips25_can_lehmann_fsm/net472 VPWR heichips25_can_lehmann_fsm/_0694_
+ VGND heichips25_can_lehmann_fsm/net1024 heichips25_can_lehmann_fsm/net365 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__3037__807 VPWR VGND net806 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2387_ VGND VPWR heichips25_can_lehmann_fsm/_0955_ heichips25_can_lehmann_fsm/net414
+ heichips25_can_lehmann_fsm/_0093_ heichips25_can_lehmann_fsm/_0659_ sg13g2_a21oi_1
XFILLER_3_118 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__3008_ net529 VGND VPWR heichips25_can_lehmann_fsm/_0233_
+ heichips25_can_lehmann_fsm__3008_/Q clknet_leaf_17_clk sg13g2_dfrbpq_1
XFILLER_47_317 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2831__545 VPWR VGND net544 sg13g2_tiehi
Xheichips25_sap3__2270_ heichips25_sap3/_1688_ heichips25_sap3/_1690_ heichips25_sap3/_1684_
+ heichips25_sap3/_1691_ VPWR VGND sg13g2_nand3_1
XFILLER_43_523 VPWR VGND sg13g2_decap_4
XFILLER_28_597 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__1985_ VPWR heichips25_sap3/_1411_ heichips25_sap3__3944_/Q VGND
+ sg13g2_inv_1
Xheichips25_sap3__3724_ heichips25_sap3/_1243_ VPWR heichips25_sap3/_0165_ VGND heichips25_sap3/_0753_
+ heichips25_sap3/_1140_ sg13g2_o21ai_1
XFILLER_3_696 VPWR VGND sg13g2_decap_4
XFILLER_2_162 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3655_ VGND VPWR heichips25_sap3/net48 heichips25_sap3/net51 heichips25_sap3/_1202_
+ heichips25_sap3/net50 sg13g2_a21oi_1
Xheichips25_sap3__2606_ heichips25_sap3/_0031_ heichips25_sap3/_0269_ heichips25_sap3/_0277_
+ heichips25_sap3/_0243_ heichips25_sap3/_1358_ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3586_ heichips25_sap3/_1111_ heichips25_sap3/_1114_ heichips25_sap3/net136
+ heichips25_sap3/_1163_ VPWR VGND heichips25_sap3/_1162_ sg13g2_nand4_1
XFILLER_47_840 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2537_ heichips25_sap3/_1883_ heichips25_sap3/_1892_ heichips25_sap3/_0213_
+ VPWR VGND sg13g2_nor2_1
XFILLER_46_350 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2468_ heichips25_sap3/_1434_ heichips25_sap3/_1782_ heichips25_sap3/_1881_
+ VPWR VGND sg13g2_and2_1
XFILLER_0_43 VPWR VGND sg13g2_decap_4
XFILLER_0_65 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2399_ heichips25_sap3/_1818_ heichips25_sap3/net77 heichips25_sap3__4025_/Q
+ heichips25_sap3/net90 heichips25_sap3__3945_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_0_98 VPWR VGND sg13g2_decap_8
XFILLER_15_770 VPWR VGND sg13g2_fill_1
XFILLER_9_63 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__4069_ heichips25_sap3__4069_/A uo_out_sap3\[0\] VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm__2310_ heichips25_can_lehmann_fsm/net327 VPWR heichips25_can_lehmann_fsm/_0619_
+ VGND heichips25_can_lehmann_fsm__2832_/Q heichips25_can_lehmann_fsm/net206 sg13g2_o21ai_1
XFILLER_30_751 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2241_ VGND VPWR heichips25_can_lehmann_fsm/net840 heichips25_can_lehmann_fsm/net170
+ heichips25_can_lehmann_fsm/_0563_ heichips25_can_lehmann_fsm/_0562_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2172_ VPWR VGND net13 heichips25_can_lehmann_fsm/_0497_
+ heichips25_can_lehmann_fsm/_0499_ heichips25_can_lehmann_fsm/net1136 heichips25_can_lehmann_fsm/_0509_
+ heichips25_can_lehmann_fsm/net175 sg13g2_a221oi_1
XFILLER_28_17 VPWR VGND sg13g2_fill_1
XFILLER_28_39 VPWR VGND sg13g2_fill_1
XFILLER_29_339 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1956_ VPWR VGND heichips25_can_lehmann_fsm/net1249 heichips25_can_lehmann_fsm/net191
+ heichips25_can_lehmann_fsm/net188 heichips25_can_lehmann_fsm/net1242 heichips25_can_lehmann_fsm/_0318_
+ heichips25_can_lehmann_fsm/net197 sg13g2_a221oi_1
XFILLER_37_372 VPWR VGND sg13g2_fill_1
XFILLER_25_523 VPWR VGND sg13g2_decap_8
XFILLER_25_534 VPWR VGND sg13g2_fill_2
Xheichips25_sap3_fanout445 heichips25_sap3/net446 heichips25_sap3/net445 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_hold1012 heichips25_sap3__4037_/Q VPWR VGND heichips25_sap3/net1011
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm__1887_ VGND VPWR heichips25_can_lehmann_fsm/_0893_ heichips25_can_lehmann_fsm/net348
+ heichips25_can_lehmann_fsm/_1200_ heichips25_can_lehmann_fsm/_0999_ sg13g2_a21oi_1
Xheichips25_sap3_fanout434 heichips25_sap3/net437 heichips25_sap3/net434 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout456 heichips25_sap3/net458 heichips25_sap3/net456 VPWR VGND
+ sg13g2_buf_1
XFILLER_12_206 VPWR VGND sg13g2_fill_1
XFILLER_25_589 VPWR VGND sg13g2_fill_1
XFILLER_21_762 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2508_ heichips25_can_lehmann_fsm/net492 VPWR heichips25_can_lehmann_fsm/_0720_
+ VGND heichips25_can_lehmann_fsm__2928_/Q heichips25_can_lehmann_fsm/net380 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2439_ VGND VPWR heichips25_can_lehmann_fsm/_0938_ heichips25_can_lehmann_fsm/net395
+ heichips25_can_lehmann_fsm/_0119_ heichips25_can_lehmann_fsm/_0685_ sg13g2_a21oi_1
XFILLER_4_438 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm_fanout382 heichips25_can_lehmann_fsm/net383 heichips25_can_lehmann_fsm/net382
+ VPWR VGND sg13g2_buf_1
XFILLER_0_600 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm_fanout371 heichips25_can_lehmann_fsm/net373 heichips25_can_lehmann_fsm/net371
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout393 heichips25_can_lehmann_fsm/net408 heichips25_can_lehmann_fsm/net393
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout360 heichips25_can_lehmann_fsm/net361 heichips25_can_lehmann_fsm/net360
+ VPWR VGND sg13g2_buf_1
Xheichips25_sap3__3440_ heichips25_sap3/net121 VPWR heichips25_sap3/_1046_ VGND heichips25_sap3/net125
+ heichips25_sap3/_1045_ sg13g2_o21ai_1
Xheichips25_sap3__3371_ VGND VPWR heichips25_sap3/net124 heichips25_sap3/_0977_ heichips25_sap3/_0980_
+ heichips25_sap3/_0979_ sg13g2_a21oi_1
XFILLER_47_169 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2322_ heichips25_sap3/_1693_ heichips25_sap3/_1736_ heichips25_sap3/_1743_
+ VPWR VGND sg13g2_and2_1
Xheichips25_sap3__2253_ heichips25_sap3/_1476_ VPWR heichips25_sap3/_1674_ VGND heichips25_sap3/net230
+ heichips25_sap3/_1496_ sg13g2_o21ai_1
XFILLER_18_83 VPWR VGND sg13g2_decap_8
XFILLER_29_895 VPWR VGND sg13g2_fill_2
XFILLER_43_342 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2883__730 VPWR VGND net729 sg13g2_tiehi
Xheichips25_sap3__2184_ heichips25_sap3/_1460_ heichips25_sap3/_1478_ heichips25_sap3/_1605_
+ VPWR VGND sg13g2_nor2_1
XFILLER_16_578 VPWR VGND sg13g2_fill_1
XFILLER_16_589 VPWR VGND sg13g2_fill_1
XFILLER_31_559 VPWR VGND sg13g2_fill_1
XFILLER_8_711 VPWR VGND sg13g2_fill_1
XFILLER_11_261 VPWR VGND sg13g2_decap_4
XFILLER_7_243 VPWR VGND sg13g2_decap_8
XFILLER_8_777 VPWR VGND sg13g2_decap_4
XFILLER_7_276 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__1968_ VPWR heichips25_sap3/_1394_ heichips25_sap3__3979_/Q VGND
+ sg13g2_inv_1
XFILLER_4_994 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3707_ heichips25_sap3/_0155_ heichips25_sap3/_1107_ heichips25_sap3/_1236_
+ heichips25_sap3/net115 heichips25_sap3/_1369_ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3638_ heichips25_sap3/_1068_ heichips25_sap3__3990_/Q heichips25_sap3/net93
+ heichips25_sap3/_0131_ VPWR VGND sg13g2_mux2_1
XFILLER_38_125 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3569_ heichips25_sap3/net119 VPWR heichips25_sap3/_1149_ VGND uio_oe_sap3\[1\]
+ heichips25_sap3/net95 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__1810_ heichips25_can_lehmann_fsm/_1126_ heichips25_can_lehmann_fsm/net294
+ heichips25_can_lehmann_fsm__2971_/Q heichips25_can_lehmann_fsm/net317 heichips25_can_lehmann_fsm__2995_/Q
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2790_ net626 VGND VPWR heichips25_can_lehmann_fsm/net1245
+ heichips25_can_lehmann_fsm__2790_/Q clknet_leaf_1_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1741_ heichips25_can_lehmann_fsm__2793_/Q heichips25_can_lehmann_fsm/_1056_
+ heichips25_can_lehmann_fsm/_1057_ heichips25_can_lehmann_fsm/_1059_ heichips25_can_lehmann_fsm/_1061_
+ VPWR VGND sg13g2_nor4_1
XFILLER_35_832 VPWR VGND sg13g2_fill_2
XFILLER_34_331 VPWR VGND sg13g2_decap_8
XFILLER_35_887 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__1672_ heichips25_can_lehmann_fsm/_0996_ heichips25_can_lehmann_fsm/net352
+ heichips25_can_lehmann_fsm/net353 VPWR VGND sg13g2_nand2_1
XFILLER_34_353 VPWR VGND sg13g2_fill_2
XFILLER_34_397 VPWR VGND sg13g2_fill_1
XFILLER_30_581 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2224_ heichips25_can_lehmann_fsm/net326 VPWR heichips25_can_lehmann_fsm/_0550_
+ VGND heichips25_can_lehmann_fsm/net1217 heichips25_can_lehmann_fsm/net161 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2155_ VGND VPWR heichips25_can_lehmann_fsm/net205 heichips25_can_lehmann_fsm/_0492_
+ heichips25_can_lehmann_fsm/_0494_ heichips25_can_lehmann_fsm/_0461_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2086_ heichips25_can_lehmann_fsm/net322 VPWR heichips25_can_lehmann_fsm/_0429_
+ VGND heichips25_can_lehmann_fsm/net345 heichips25_can_lehmann_fsm/net179 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2988_ net672 VGND VPWR heichips25_can_lehmann_fsm/_0213_
+ heichips25_can_lehmann_fsm__2988_/Q clknet_leaf_18_clk sg13g2_dfrbpq_1
Xheichips25_sap3_fanout220 heichips25_sap3/_1642_ heichips25_sap3/net220 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout231 heichips25_sap3/net233 heichips25_sap3/net231 VPWR VGND
+ sg13g2_buf_1
Xheichips25_can_lehmann_fsm__1939_ heichips25_can_lehmann_fsm/_1090_ VPWR heichips25_can_lehmann_fsm/_0302_
+ VGND heichips25_can_lehmann_fsm/net219 heichips25_can_lehmann_fsm/_0301_ sg13g2_o21ai_1
Xheichips25_sap3_fanout242 heichips25_sap3/_1520_ heichips25_sap3/net242 VPWR VGND
+ sg13g2_buf_1
XFILLER_13_515 VPWR VGND sg13g2_decap_8
Xheichips25_sap3_fanout264 heichips25_sap3__3926_/Q heichips25_sap3/net264 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout253 heichips25_sap3__4063_/Q heichips25_sap3/net253 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout275 heichips25_sap3__3906_/Q heichips25_sap3/net275 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout286 heichips25_sap3__3900_/Q heichips25_sap3/net286 VPWR VGND
+ sg13g2_buf_1
Xrebuffer830 uio_oe_sap3\[5\] net829 VPWR VGND sg13g2_buf_2
XFILLER_5_714 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2940_ heichips25_sap3/_0579_ heichips25_sap3/_0576_ heichips25_sap3/_0578_
+ VPWR VGND sg13g2_xnor2_1
Xheichips25_sap3__2871_ heichips25_sap3/_0511_ heichips25_sap3/_0512_ heichips25_sap3/_0507_
+ heichips25_sap3/_0513_ VPWR VGND sg13g2_nand3_1
XFILLER_5_769 VPWR VGND sg13g2_decap_8
Xclkbuf_5_17__f_heichips25_sap3\_sap_3_inst.alu_inst.clk heichips25_sap3__3922_/CLK
+ clknet_4_8_0_heichips25_sap3\/sap_3_inst.alu_inst.clk VPWR VGND sg13g2_buf_16
Xheichips25_can_lehmann_fsm_fanout190 heichips25_can_lehmann_fsm/_0307_ heichips25_can_lehmann_fsm/net190
+ VPWR VGND sg13g2_buf_1
XFILLER_0_463 VPWR VGND sg13g2_fill_1
XFILLER_1_975 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3423_ heichips25_sap3/_0078_ heichips25_sap3/_1023_ heichips25_sap3/_1029_
+ heichips25_sap3/_0748_ heichips25_sap3/_1412_ VPWR VGND sg13g2_a22oi_1
XFILLER_49_979 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3354_ heichips25_sap3/_0961_ heichips25_sap3/_0962_ heichips25_sap3/_0960_
+ heichips25_sap3/_0963_ VPWR VGND sg13g2_nand3_1
Xheichips25_sap3__2305_ heichips25_sap3/net264 heichips25_sap3/_1725_ heichips25_sap3/_1726_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__3285_ VPWR VGND heichips25_sap3__3988_/Q heichips25_sap3/_0896_
+ heichips25_sap3/net133 heichips25_sap3__3980_/Q heichips25_sap3/_0897_ heichips25_sap3/net141
+ sg13g2_a221oi_1
Xheichips25_sap3__2236_ VGND VPWR heichips25_sap3/net238 heichips25_sap3/_1656_ heichips25_sap3/_1657_
+ heichips25_sap3/_1641_ sg13g2_a21oi_1
Xheichips25_sap3__2167_ heichips25_sap3/_1571_ heichips25_sap3/_1584_ heichips25_sap3/_1587_
+ heichips25_sap3/_1588_ VPWR VGND sg13g2_nor3_1
XFILLER_32_835 VPWR VGND sg13g2_fill_1
XFILLER_31_345 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2098_ heichips25_sap3/_1515_ heichips25_sap3/_1517_ heichips25_sap3/_1519_
+ VPWR VGND sg13g2_nor2_1
XFILLER_12_581 VPWR VGND sg13g2_fill_1
XFILLER_6_97 VPWR VGND sg13g2_decap_8
XFILLER_39_434 VPWR VGND sg13g2_fill_1
XFILLER_39_423 VPWR VGND sg13g2_decap_8
XFILLER_6_1024 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2911_ net673 VGND VPWR heichips25_can_lehmann_fsm/net967
+ heichips25_can_lehmann_fsm__2911_/Q clknet_leaf_15_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2842_ net811 VGND VPWR heichips25_can_lehmann_fsm/_0067_
+ heichips25_can_lehmann_fsm__2842_/Q clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_13_0 VPWR VGND sg13g2_fill_2
XFILLER_26_106 VPWR VGND sg13g2_fill_1
XFILLER_26_128 VPWR VGND sg13g2_decap_8
XFILLER_27_629 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2773_ uo_out_fsm\[1\] heichips25_can_lehmann_fsm/net321
+ heichips25_can_lehmann_fsm/_0287_ VPWR VGND sg13g2_and2_1
Xheichips25_can_lehmann_fsm__1724_ heichips25_can_lehmann_fsm/net1181 heichips25_can_lehmann_fsm__2822_/Q
+ heichips25_can_lehmann_fsm/_1044_ heichips25_can_lehmann_fsm/_1045_ VPWR VGND sg13g2_nor3_1
XFILLER_23_802 VPWR VGND sg13g2_fill_1
XFILLER_34_161 VPWR VGND sg13g2_fill_2
XFILLER_23_835 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__1655_ VPWR heichips25_can_lehmann_fsm/_0979_ heichips25_can_lehmann_fsm__2791_/Q
+ VGND sg13g2_inv_1
XFILLER_22_345 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__1586_ VPWR heichips25_can_lehmann_fsm/_0910_ heichips25_can_lehmann_fsm/net1060
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__2207_ VGND VPWR heichips25_can_lehmann_fsm/net161 heichips25_can_lehmann_fsm/_0535_
+ heichips25_can_lehmann_fsm/_0036_ heichips25_can_lehmann_fsm/_0536_ sg13g2_a21oi_1
XFILLER_1_205 VPWR VGND sg13g2_decap_8
XFILLER_9_8 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2138_ heichips25_can_lehmann_fsm/_0477_ heichips25_can_lehmann_fsm/net349
+ heichips25_can_lehmann_fsm__2980_/Q VPWR VGND sg13g2_nand2b_1
Xheichips25_can_lehmann_fsm__2069_ VPWR VGND heichips25_can_lehmann_fsm/net346 heichips25_can_lehmann_fsm/net182
+ heichips25_can_lehmann_fsm/net190 heichips25_can_lehmann_fsm/net1255 heichips25_can_lehmann_fsm/_0415_
+ heichips25_can_lehmann_fsm/net199 sg13g2_a221oi_1
XFILLER_17_139 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3070_ heichips25_sap3/_1365_ heichips25_sap3/_1480_ heichips25_sap3/_1619_
+ heichips25_sap3/_0683_ VPWR VGND sg13g2_nor3_1
XFILLER_26_651 VPWR VGND sg13g2_fill_2
XFILLER_26_673 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2021_ heichips25_sap3/_1442_ heichips25_sap3/net263 heichips25_sap3/net261
+ VPWR VGND sg13g2_nand2_1
XFILLER_13_301 VPWR VGND sg13g2_decap_4
XFILLER_25_161 VPWR VGND sg13g2_fill_1
XFILLER_40_142 VPWR VGND sg13g2_fill_1
XFILLER_40_120 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm_hold1151 heichips25_can_lehmann_fsm__3008_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1150 sg13g2_dlygate4sd3_1
XFILLER_15_51 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm_hold1140 heichips25_can_lehmann_fsm__3007_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1139 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1184 heichips25_can_lehmann_fsm__2854_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1183 sg13g2_dlygate4sd3_1
XFILLER_40_175 VPWR VGND sg13g2_decap_8
XFILLER_40_164 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_hold1173 heichips25_can_lehmann_fsm__3035_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1172 sg13g2_dlygate4sd3_1
XFILLER_13_389 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm_hold1162 heichips25_can_lehmann_fsm/_0259_ VPWR VGND heichips25_can_lehmann_fsm/net1161
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1195 heichips25_can_lehmann_fsm__2824_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1194 sg13g2_dlygate4sd3_1
Xheichips25_sap3__3972_ heichips25_sap3/net443 VGND VPWR heichips25_sap3/_0113_ heichips25_sap3__3972_/Q
+ heichips25_sap3__3988_/CLK sg13g2_dfrbpq_1
Xheichips25_sap3_hold893 heichips25_sap3/_0177_ VPWR VGND heichips25_sap3/net892 sg13g2_dlygate4sd3_1
Xheichips25_sap3__2923_ VPWR heichips25_sap3/_0562_ heichips25_sap3/_0561_ VGND sg13g2_inv_1
Xheichips25_sap3_fanout81 heichips25_sap3/net82 heichips25_sap3/net81 VPWR VGND sg13g2_buf_1
XFILLER_5_577 VPWR VGND sg13g2_fill_1
Xheichips25_sap3_fanout70 heichips25_sap3/_0440_ heichips25_sap3/net70 VPWR VGND sg13g2_buf_1
Xheichips25_sap3__2854_ heichips25_sap3/net70 heichips25_sap3/net285 heichips25_sap3/_0496_
+ heichips25_sap3/_0042_ VPWR VGND sg13g2_a21o_1
Xheichips25_sap3__2785_ heichips25_sap3/net238 heichips25_sap3/_1643_ heichips25_sap3/_1449_
+ heichips25_sap3/_0430_ VPWR VGND sg13g2_nand3_1
Xheichips25_sap3_fanout92 heichips25_sap3/_1733_ heichips25_sap3/net92 VPWR VGND sg13g2_buf_1
XFILLER_0_260 VPWR VGND sg13g2_decap_8
XFILLER_48_231 VPWR VGND sg13g2_fill_1
XFILLER_49_798 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3406_ VPWR VGND heichips25_sap3__3961_/Q heichips25_sap3/_1012_
+ heichips25_sap3/_0760_ heichips25_sap3__3953_/Q heichips25_sap3/_1013_ heichips25_sap3/net110
+ sg13g2_a221oi_1
XFILLER_36_459 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3337_ heichips25_sap3/_0947_ heichips25_sap3/_0819_ heichips25_sap3/_0934_
+ VPWR VGND sg13g2_xnor2_1
Xheichips25_sap3__3268_ heichips25_sap3/_0881_ heichips25_sap3/_0715_ heichips25_sap3/_0880_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__2219_ heichips25_sap3/_1450_ VPWR heichips25_sap3/_1640_ VGND heichips25_sap3/_1501_
+ heichips25_sap3/_1506_ sg13g2_o21ai_1
XFILLER_17_684 VPWR VGND sg13g2_fill_1
XFILLER_32_632 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3199_ heichips25_sap3/_0717_ heichips25_sap3/net151 heichips25_sap3__4022_/Q
+ heichips25_sap3/_0812_ VPWR VGND sg13g2_nand3_1
XFILLER_9_894 VPWR VGND sg13g2_decap_8
XFILLER_8_393 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__3041_ net742 VGND VPWR heichips25_can_lehmann_fsm/_0266_
+ heichips25_can_lehmann_fsm__3041_/Q clknet_leaf_22_clk sg13g2_dfrbpq_1
XFILLER_28_1014 VPWR VGND sg13g2_fill_1
XFILLER_39_253 VPWR VGND sg13g2_decap_8
XFILLER_36_17 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2825_ net556 VGND VPWR heichips25_can_lehmann_fsm/_0050_
+ heichips25_can_lehmann_fsm__2825_/Q clknet_leaf_10_clk sg13g2_dfrbpq_1
XFILLER_27_448 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2756_ heichips25_can_lehmann_fsm/net498 VPWR heichips25_can_lehmann_fsm/_0844_
+ VGND heichips25_can_lehmann_fsm__3052_/Q heichips25_can_lehmann_fsm/net384 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__1707_ VGND VPWR heichips25_can_lehmann_fsm/_1031_ heichips25_can_lehmann_fsm/_1029_
+ heichips25_can_lehmann_fsm/_1016_ sg13g2_or2_1
Xheichips25_can_lehmann_fsm__2687_ VGND VPWR heichips25_can_lehmann_fsm/_0874_ heichips25_can_lehmann_fsm/net398
+ heichips25_can_lehmann_fsm/_0243_ heichips25_can_lehmann_fsm/_0809_ sg13g2_a21oi_1
XFILLER_22_142 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1638_ VPWR heichips25_can_lehmann_fsm/_0962_ heichips25_can_lehmann_fsm/net898
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__1569_ VPWR heichips25_can_lehmann_fsm/_0893_ heichips25_can_lehmann_fsm/net985
+ VGND sg13g2_inv_1
XFILLER_2_514 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2570_ VGND VPWR heichips25_sap3/net215 heichips25_sap3/net45 heichips25_sap3/_0244_
+ heichips25_sap3/_0243_ sg13g2_a21oi_1
Xheichips25_sap3__3122_ VGND VPWR heichips25_sap3/_0735_ heichips25_sap3/_1635_ heichips25_sap3/_1532_
+ sg13g2_or2_1
XFILLER_26_470 VPWR VGND sg13g2_fill_1
XFILLER_26_492 VPWR VGND sg13g2_decap_8
XFILLER_42_952 VPWR VGND sg13g2_fill_1
XFILLER_13_142 VPWR VGND sg13g2_fill_2
XFILLER_14_654 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3053_ VGND VPWR heichips25_sap3/net241 heichips25_sap3/_0659_ heichips25_sap3/_0666_
+ heichips25_sap3/_0664_ sg13g2_a21oi_1
XFILLER_41_484 VPWR VGND sg13g2_decap_4
XFILLER_13_175 VPWR VGND sg13g2_fill_1
XFILLER_14_687 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2004_ VPWR heichips25_sap3/_1429_ heichips25_sap3__4074_/A VGND
+ sg13g2_inv_1
XFILLER_42_82 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3955_ heichips25_sap3/net456 VGND VPWR heichips25_sap3/_0096_ heichips25_sap3__3955_/Q
+ clkload28/A sg13g2_dfrbpq_1
Xheichips25_sap3__3886_ heichips25_sap3/net453 VGND VPWR heichips25_sap3/_0027_ heichips25_sap3__3886_/Q
+ clkload25/A sg13g2_dfrbpq_1
Xheichips25_sap3__2906_ heichips25_sap3/_0545_ VPWR heichips25_sap3/_0546_ VGND heichips25_sap3/_0379_
+ heichips25_sap3/_0522_ sg13g2_o21ai_1
Xheichips25_sap3__2837_ heichips25_sap3/_0480_ heichips25_sap3/_0361_ heichips25_sap3/_0445_
+ VPWR VGND sg13g2_nand2_1
X_23__509 VPWR VGND net508 sg13g2_tielo
XFILLER_3_21 VPWR VGND sg13g2_decap_8
XFILLER_3_65 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2768_ VGND VPWR heichips25_sap3/_1374_ heichips25_sap3__3922_/Q
+ heichips25_sap3/_0414_ heichips25_sap3/_0411_ sg13g2_a21oi_1
Xheichips25_sap3__2699_ heichips25_sap3/_0345_ heichips25_sap3/_1888_ heichips25_sap3/_0344_
+ VPWR VGND sg13g2_nand2_1
Xclkbuf_5_0__f_heichips25_sap3\_sap_3_inst.alu_inst.clk heichips25_sap3__4013_/CLK
+ clknet_4_0_0_heichips25_sap3\/sap_3_inst.alu_inst.clk VPWR VGND sg13g2_buf_16
XFILLER_49_584 VPWR VGND sg13g2_fill_2
XFILLER_49_562 VPWR VGND sg13g2_decap_8
XFILLER_3_1005 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2610_ heichips25_can_lehmann_fsm/net485 VPWR heichips25_can_lehmann_fsm/_0771_
+ VGND heichips25_can_lehmann_fsm__2980_/Q heichips25_can_lehmann_fsm/net413 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2541_ VGND VPWR heichips25_can_lehmann_fsm/_0912_ heichips25_can_lehmann_fsm/net356
+ heichips25_can_lehmann_fsm/_0170_ heichips25_can_lehmann_fsm/_0736_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2472_ heichips25_can_lehmann_fsm/net488 VPWR heichips25_can_lehmann_fsm/_0702_
+ VGND heichips25_can_lehmann_fsm__2910_/Q heichips25_can_lehmann_fsm/net377 sg13g2_o21ai_1
XFILLER_20_635 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__3024_ net690 VGND VPWR heichips25_can_lehmann_fsm/_0249_
+ heichips25_can_lehmann_fsm__3024_/Q clknet_leaf_7_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2808_ net590 VGND VPWR heichips25_can_lehmann_fsm/net1193
+ heichips25_can_lehmann_fsm__2808_/Q clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_43_716 VPWR VGND sg13g2_fill_1
XFILLER_43_705 VPWR VGND sg13g2_decap_8
XFILLER_15_407 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__2944__560 VPWR VGND net559 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2739_ VGND VPWR heichips25_can_lehmann_fsm/_0860_ heichips25_can_lehmann_fsm/net355
+ heichips25_can_lehmann_fsm/_0269_ heichips25_can_lehmann_fsm/_0835_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2842__812 VPWR VGND net811 sg13g2_tiehi
Xheichips25_can_lehmann_fsm_hold867 heichips25_can_lehmann_fsm/_0120_ VPWR VGND heichips25_can_lehmann_fsm/net866
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold856 heichips25_can_lehmann_fsm__2997_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net855 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold845 heichips25_can_lehmann_fsm__2999_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net844 sg13g2_dlygate4sd3_1
XFILLER_10_156 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_hold878 heichips25_can_lehmann_fsm__3042_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net877 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold889 heichips25_can_lehmann_fsm/_0195_ VPWR VGND heichips25_can_lehmann_fsm/net888
+ sg13g2_dlygate4sd3_1
Xheichips25_sap3__3740_ VGND VPWR heichips25_sap3/net1176 heichips25_sap3/_1246_ heichips25_sap3/_0170_
+ heichips25_sap3/_1254_ sg13g2_a21oi_1
Xheichips25_sap3__3671_ heichips25_sap3/_1212_ heichips25_sap3/_1214_ heichips25_sap3/_1215_
+ VPWR VGND sg13g2_and2_1
XFILLER_2_333 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2622_ VGND VPWR heichips25_sap3/net1130 heichips25_sap3/_1431_ heichips25_sap3/_0291_
+ heichips25_sap3/_0290_ sg13g2_a21oi_1
Xheichips25_sap3__2553_ heichips25_sap3/_0228_ heichips25_sap3/net82 heichips25_sap3__3966_/Q
+ heichips25_sap3/net83 heichips25_sap3__3958_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2484_ heichips25_sap3/_1893_ VPWR heichips25_sap3/_1897_ VGND heichips25_sap3/net159
+ heichips25_sap3/_1896_ sg13g2_o21ai_1
XFILLER_19_735 VPWR VGND sg13g2_fill_1
XFILLER_37_71 VPWR VGND sg13g2_decap_8
XFILLER_18_267 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3105_ heichips25_sap3/_0718_ heichips25_sap3/_0697_ heichips25_sap3/_0714_
+ heichips25_sap3/_0716_ VPWR VGND sg13g2_and3_1
XFILLER_18_1013 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3036_ heichips25_sap3/_0649_ heichips25_sap3/_1580_ heichips25_sap3/_1486_
+ heichips25_sap3/_1532_ heichips25_sap3/_1513_ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2923__644 VPWR VGND net643 sg13g2_tiehi
Xheichips25_sap3__3938_ heichips25_sap3/net440 VGND VPWR heichips25_sap3/_0079_ heichips25_sap3__3938_/Q
+ heichips25_sap3__4018_/CLK sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2893__710 VPWR VGND net709 sg13g2_tiehi
XFILLER_5_182 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3869_ heichips25_sap3__3888_/Q heichips25_sap3/net1105 heichips25_sap3/net341
+ heichips25_sap3/_0196_ VPWR VGND sg13g2_mux2_1
XFILLER_38_2 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1972_ heichips25_can_lehmann_fsm/net322 VPWR heichips25_can_lehmann_fsm/_0332_
+ VGND heichips25_can_lehmann_fsm/net1260 heichips25_can_lehmann_fsm/net178 sg13g2_o21ai_1
XFILLER_37_587 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2524_ heichips25_can_lehmann_fsm/net483 VPWR heichips25_can_lehmann_fsm/_0728_
+ VGND heichips25_can_lehmann_fsm/net1079 heichips25_can_lehmann_fsm/net375 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2455_ VGND VPWR heichips25_can_lehmann_fsm/_0934_ heichips25_can_lehmann_fsm/net404
+ heichips25_can_lehmann_fsm/_0127_ heichips25_can_lehmann_fsm/_0693_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2386_ heichips25_can_lehmann_fsm/net480 VPWR heichips25_can_lehmann_fsm/_0659_
+ VGND heichips25_can_lehmann_fsm/net1068 heichips25_can_lehmann_fsm/net414 sg13g2_o21ai_1
XFILLER_20_498 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__3007_ net537 VGND VPWR heichips25_can_lehmann_fsm/net1140
+ heichips25_can_lehmann_fsm__3007_/Q clknet_leaf_15_clk sg13g2_dfrbpq_1
XFILLER_28_554 VPWR VGND sg13g2_decap_4
XFILLER_12_911 VPWR VGND sg13g2_fill_1
XFILLER_12_944 VPWR VGND sg13g2_decap_8
XFILLER_7_458 VPWR VGND sg13g2_decap_4
XFILLER_7_447 VPWR VGND sg13g2_fill_2
XFILLER_8_959 VPWR VGND sg13g2_decap_4
XFILLER_23_84 VPWR VGND sg13g2_fill_1
XFILLER_7_469 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__1984_ VPWR heichips25_sap3/_1410_ heichips25_sap3__3952_/Q VGND
+ sg13g2_inv_1
XFILLER_48_1028 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3723_ heichips25_sap3/_1243_ heichips25_sap3__4024_/Q heichips25_sap3/_0753_
+ VPWR VGND sg13g2_nand2_1
XFILLER_3_664 VPWR VGND sg13g2_fill_1
XFILLER_3_631 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3654_ heichips25_sap3/_0137_ heichips25_sap3/_1095_ heichips25_sap3/_1201_
+ heichips25_sap3/net112 heichips25_sap3/_1387_ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2605_ VGND VPWR heichips25_sap3/_1802_ heichips25_sap3/_0276_ heichips25_sap3/_0277_
+ heichips25_sap3/_0243_ sg13g2_a21oi_1
Xheichips25_sap3__3585_ heichips25_sap3/_1161_ VPWR heichips25_sap3/_1162_ VGND uio_oe_sap3\[4\]
+ heichips25_sap3/net95 sg13g2_o21ai_1
XFILLER_38_329 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2536_ VPWR heichips25_sap3/_0212_ uio_out_sap3\[0\] VGND sg13g2_inv_1
XFILLER_47_863 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2467_ heichips25_sap3__3928_/Q heichips25_sap3/_1879_ heichips25_sap3/_1880_
+ VPWR VGND sg13g2_and2_1
XFILLER_0_22 VPWR VGND sg13g2_decap_8
XFILLER_46_384 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2398_ heichips25_sap3/_1817_ heichips25_sap3/net75 heichips25_sap3__3993_/Q
+ heichips25_sap3/net84 heichips25_sap3__3969_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_14_270 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3019_ VGND VPWR heichips25_sap3/_1364_ heichips25_sap3/net232 heichips25_sap3/_0068_
+ heichips25_sap3/_0635_ sg13g2_a21oi_1
XFILLER_30_774 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2240_ heichips25_can_lehmann_fsm/net170 heichips25_can_lehmann_fsm/_0561_
+ heichips25_can_lehmann_fsm/_0562_ VPWR VGND sg13g2_nor2_1
Xheichips25_can_lehmann_fsm__2171_ heichips25_can_lehmann_fsm/_0508_ heichips25_can_lehmann_fsm/net164
+ heichips25_can_lehmann_fsm/_0507_ VPWR VGND sg13g2_nand2_1
X_29__515 VPWR VGND net514 sg13g2_tielo
XFILLER_29_318 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1955_ heichips25_can_lehmann_fsm/_0317_ heichips25_can_lehmann_fsm/net184
+ heichips25_can_lehmann_fsm/_0316_ VPWR VGND sg13g2_nand2_1
Xheichips25_can_lehmann_fsm__1886_ heichips25_can_lehmann_fsm/_1199_ heichips25_can_lehmann_fsm/_0941_
+ heichips25_can_lehmann_fsm/net302 VPWR VGND sg13g2_nand2_1
Xheichips25_sap3_fanout446 _01_ heichips25_sap3/net446 VPWR VGND sg13g2_buf_1
Xheichips25_sap3_hold1013 heichips25_sap3/_0178_ VPWR VGND heichips25_sap3/net1012
+ sg13g2_dlygate4sd3_1
XFILLER_44_39 VPWR VGND sg13g2_fill_2
Xheichips25_sap3_fanout435 heichips25_sap3/net437 heichips25_sap3/net435 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout457 heichips25_sap3/net458 heichips25_sap3/net457 VPWR VGND
+ sg13g2_buf_1
Xheichips25_can_lehmann_fsm__2507_ VGND VPWR heichips25_can_lehmann_fsm/_0921_ heichips25_can_lehmann_fsm/net421
+ heichips25_can_lehmann_fsm/_0153_ heichips25_can_lehmann_fsm/_0719_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2438_ heichips25_can_lehmann_fsm/net464 VPWR heichips25_can_lehmann_fsm/_0685_
+ VGND heichips25_can_lehmann_fsm__2894_/Q heichips25_can_lehmann_fsm/net394 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2369_ VGND VPWR heichips25_can_lehmann_fsm/_0959_ heichips25_can_lehmann_fsm/net388
+ heichips25_can_lehmann_fsm/_0084_ heichips25_can_lehmann_fsm/_0650_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm_fanout350 heichips25_can_lehmann_fsm__2777_/Q heichips25_can_lehmann_fsm/net350
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout383 heichips25_can_lehmann_fsm/net388 heichips25_can_lehmann_fsm/net383
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout372 heichips25_can_lehmann_fsm/net373 heichips25_can_lehmann_fsm/net372
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout361 heichips25_can_lehmann_fsm/net362 heichips25_can_lehmann_fsm/net361
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout394 heichips25_can_lehmann_fsm/net397 heichips25_can_lehmann_fsm/net394
+ VPWR VGND sg13g2_buf_1
Xheichips25_sap3__3370_ heichips25_sap3/net121 VPWR heichips25_sap3/_0979_ VGND heichips25_sap3/net124
+ heichips25_sap3/_0978_ sg13g2_o21ai_1
Xheichips25_sap3__2321_ heichips25_sap3/_1712_ heichips25_sap3/_1731_ heichips25_sap3/_1693_
+ heichips25_sap3/_1742_ VPWR VGND sg13g2_nand3_1
Xheichips25_sap3__2252_ heichips25_sap3/_1666_ heichips25_sap3/_1669_ heichips25_sap3/_1663_
+ heichips25_sap3/_1673_ VPWR VGND heichips25_sap3/_1672_ sg13g2_nand4_1
XFILLER_28_362 VPWR VGND sg13g2_fill_2
XFILLER_16_546 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2183_ VGND VPWR heichips25_sap3/net243 heichips25_sap3/_1603_ heichips25_sap3/_1604_
+ heichips25_sap3/_1577_ sg13g2_a21oi_1
XFILLER_31_516 VPWR VGND sg13g2_decap_4
XFILLER_31_538 VPWR VGND sg13g2_decap_8
XFILLER_34_50 VPWR VGND sg13g2_decap_4
XFILLER_7_233 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__1967_ VPWR heichips25_sap3/_1393_ heichips25_sap3__4019_/Q VGND
+ sg13g2_inv_1
Xheichips25_sap3__3706_ uio_oe_sap3\[3\] heichips25_sap3/net115 heichips25_sap3/_1236_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__3637_ VGND VPWR heichips25_sap3/_0888_ heichips25_sap3/_1159_ heichips25_sap3/_1191_
+ heichips25_sap3/_1068_ sg13g2_a21oi_1
XFILLER_15_4 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3568_ heichips25_sap3/_1142_ VPWR heichips25_sap3/_0104_ VGND heichips25_sap3/_1143_
+ heichips25_sap3/_1148_ sg13g2_o21ai_1
Xheichips25_sap3__2519_ heichips25_sap3/_1928_ heichips25_sap3/_1929_ heichips25_sap3/_1930_
+ VPWR VGND sg13g2_and2_1
Xheichips25_can_lehmann_fsm__1740_ heichips25_can_lehmann_fsm/_1058_ heichips25_can_lehmann_fsm/_1059_
+ heichips25_can_lehmann_fsm/_1060_ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__3499_ heichips25_sap3/_1093_ heichips25_sap3/_1094_ heichips25_sap3/_1095_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_can_lehmann_fsm__1671_ heichips25_can_lehmann_fsm/net351 heichips25_can_lehmann_fsm/net348
+ heichips25_can_lehmann_fsm/_0995_ VPWR VGND heichips25_can_lehmann_fsm/net353 sg13g2_nand3b_1
XFILLER_22_549 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2223_ heichips25_can_lehmann_fsm/_0549_ heichips25_can_lehmann_fsm/net165
+ heichips25_can_lehmann_fsm/_0548_ heichips25_can_lehmann_fsm/net176 heichips25_can_lehmann_fsm/net1050
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2154_ heichips25_can_lehmann_fsm/_0493_ heichips25_can_lehmann_fsm/net205
+ heichips25_can_lehmann_fsm/_0492_ VPWR VGND sg13g2_xnor2_1
Xheichips25_can_lehmann_fsm__2085_ heichips25_can_lehmann_fsm/_0428_ heichips25_can_lehmann_fsm/net186
+ heichips25_can_lehmann_fsm/_0427_ heichips25_can_lehmann_fsm/net199 heichips25_can_lehmann_fsm/net1266
+ VPWR VGND sg13g2_a22oi_1
XFILLER_39_28 VPWR VGND sg13g2_fill_2
XFILLER_29_104 VPWR VGND sg13g2_fill_2
XFILLER_29_115 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2987_ net676 VGND VPWR heichips25_can_lehmann_fsm/net890
+ heichips25_can_lehmann_fsm__2987_/Q clknet_leaf_17_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__1938_ VGND VPWR heichips25_can_lehmann_fsm/_0945_ heichips25_can_lehmann_fsm/net302
+ heichips25_can_lehmann_fsm/_0301_ heichips25_can_lehmann_fsm/_0300_ sg13g2_a21oi_1
Xheichips25_sap3_fanout221 heichips25_sap3/_1642_ heichips25_sap3/net221 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout232 heichips25_sap3/net233 heichips25_sap3/net232 VPWR VGND
+ sg13g2_buf_1
XFILLER_41_814 VPWR VGND sg13g2_decap_8
Xheichips25_sap3_fanout254 heichips25_sap3__3893_/Q heichips25_sap3/net254 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout243 heichips25_sap3/_1512_ heichips25_sap3/net243 VPWR VGND
+ sg13g2_buf_2
Xheichips25_sap3_fanout265 heichips25_sap3__3926_/Q heichips25_sap3/net265 VPWR VGND
+ sg13g2_buf_1
Xheichips25_can_lehmann_fsm__1869_ heichips25_can_lehmann_fsm/_0999_ heichips25_can_lehmann_fsm/_1163_
+ heichips25_can_lehmann_fsm/_0996_ heichips25_can_lehmann_fsm/_1184_ VPWR VGND sg13g2_nand3_1
XFILLER_26_899 VPWR VGND sg13g2_fill_1
Xheichips25_sap3_fanout276 heichips25_sap3__3905_/Q heichips25_sap3/net276 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout287 heichips25_sap3__3900_/Q heichips25_sap3/net287 VPWR VGND
+ sg13g2_buf_1
Xheichips25_can_lehmann_fsm__2800__607 VPWR VGND net606 sg13g2_tiehi
Xheichips25_sap3__2870_ heichips25_sap3/_0512_ heichips25_sap3/_0442_ heichips25_sap3/_1367_
+ heichips25_sap3/_0416_ heichips25_sap3/net280 VPWR VGND sg13g2_a22oi_1
XFILLER_4_203 VPWR VGND sg13g2_decap_8
XFILLER_1_954 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm_fanout180 heichips25_can_lehmann_fsm/_0313_ heichips25_can_lehmann_fsm/net180
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout191 heichips25_can_lehmann_fsm/net192 heichips25_can_lehmann_fsm/net191
+ VPWR VGND sg13g2_buf_1
Xheichips25_sap3__3422_ heichips25_sap3/_0748_ heichips25_sap3/_1027_ heichips25_sap3/_1028_
+ heichips25_sap3/_1029_ VPWR VGND sg13g2_nor3_1
XFILLER_49_969 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2850__796 VPWR VGND net795 sg13g2_tiehi
Xheichips25_sap3__3353_ heichips25_sap3/_0962_ heichips25_sap3/net135 heichips25_sap3__3967_/Q
+ heichips25_sap3/net139 heichips25_sap3__3975_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_29_72 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2304_ heichips25_sap3/net245 heichips25_sap3/_1551_ heichips25_sap3/_1463_
+ heichips25_sap3/_1725_ VPWR VGND sg13g2_nand3_1
Xheichips25_sap3__3284_ heichips25_sap3/_0892_ VPWR heichips25_sap3/_0896_ VGND heichips25_sap3/_1386_
+ heichips25_sap3/net115 sg13g2_o21ai_1
XFILLER_44_652 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2235_ VPWR heichips25_sap3/_1656_ heichips25_sap3/_1655_ VGND sg13g2_inv_1
XFILLER_43_195 VPWR VGND sg13g2_fill_2
XFILLER_43_173 VPWR VGND sg13g2_fill_1
XFILLER_43_162 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2166_ heichips25_sap3/_1585_ heichips25_sap3/_1586_ heichips25_sap3/_1579_
+ heichips25_sap3/_1587_ VPWR VGND sg13g2_nand3_1
XFILLER_31_302 VPWR VGND sg13g2_decap_8
XFILLER_31_324 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2097_ VGND VPWR heichips25_sap3/_1518_ heichips25_sap3/_1511_ heichips25_sap3/_1506_
+ sg13g2_or2_1
XFILLER_8_531 VPWR VGND sg13g2_decap_8
XFILLER_6_65 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2999_ heichips25_sap3/_0626_ VPWR heichips25_sap3/_0057_ VGND heichips25_sap3/_1396_
+ heichips25_sap3/net201 sg13g2_o21ai_1
XFILLER_3_280 VPWR VGND sg13g2_decap_8
XFILLER_6_1014 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2910_ net675 VGND VPWR heichips25_can_lehmann_fsm/net910
+ heichips25_can_lehmann_fsm__2910_/Q clknet_leaf_15_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2841_ net813 VGND VPWR heichips25_can_lehmann_fsm/net1089
+ heichips25_can_lehmann_fsm__2841_/Q clknet_leaf_4_clk sg13g2_dfrbpq_1
Xheichips25_can_lehmann_fsm__2772_ uo_out_fsm\[0\] heichips25_can_lehmann_fsm/net321
+ heichips25_can_lehmann_fsm/_0286_ VPWR VGND sg13g2_and2_1
Xheichips25_can_lehmann_fsm__1723_ heichips25_can_lehmann_fsm__2821_/Q heichips25_can_lehmann_fsm__2820_/Q
+ heichips25_can_lehmann_fsm__2819_/Q heichips25_can_lehmann_fsm__2818_/Q heichips25_can_lehmann_fsm/_1044_
+ VPWR VGND sg13g2_or4_1
Xheichips25_can_lehmann_fsm__1654_ VPWR heichips25_can_lehmann_fsm/_0978_ heichips25_can_lehmann_fsm__2792_/Q
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__1585_ VPWR heichips25_can_lehmann_fsm/_0909_ heichips25_can_lehmann_fsm/net1077
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__2206_ heichips25_can_lehmann_fsm/net325 VPWR heichips25_can_lehmann_fsm/_0536_
+ VGND heichips25_can_lehmann_fsm/net1180 heichips25_can_lehmann_fsm/net161 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2137_ heichips25_can_lehmann_fsm/_0475_ heichips25_can_lehmann_fsm/_1138_
+ heichips25_can_lehmann_fsm/_0468_ heichips25_can_lehmann_fsm/_0476_ VPWR VGND sg13g2_a21o_1
Xheichips25_can_lehmann_fsm__2068_ heichips25_can_lehmann_fsm/_0414_ heichips25_can_lehmann_fsm/net186
+ heichips25_can_lehmann_fsm/_0402_ heichips25_can_lehmann_fsm/net195 net12 VPWR VGND
+ sg13g2_a22oi_1
XFILLER_38_490 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2020_ heichips25_sap3/net262 heichips25_sap3/net261 heichips25_sap3/_1441_
+ VPWR VGND sg13g2_and2_1
XFILLER_26_685 VPWR VGND sg13g2_decap_8
XFILLER_41_666 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_hold1130 heichips25_can_lehmann_fsm__3013_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1129 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1141 heichips25_can_lehmann_fsm/_0232_ VPWR VGND heichips25_can_lehmann_fsm/net1140
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1174 heichips25_can_lehmann_fsm__2821_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1173 sg13g2_dlygate4sd3_1
XFILLER_15_85 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm_hold1152 heichips25_can_lehmann_fsm__3046_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1151 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1185 heichips25_can_lehmann_fsm/_0576_ VPWR VGND heichips25_can_lehmann_fsm/net1184
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1196 heichips25_can_lehmann_fsm__2820_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1195 sg13g2_dlygate4sd3_1
Xheichips25_sap3__3971_ heichips25_sap3/net456 VGND VPWR heichips25_sap3/_0112_ heichips25_sap3__3971_/Q
+ heichips25_sap3__3990_/CLK sg13g2_dfrbpq_1
Xheichips25_sap3__2922_ heichips25_sap3/_0369_ heichips25_sap3/_0350_ heichips25_sap3/_0561_
+ VPWR VGND sg13g2_xor2_1
XFILLER_5_523 VPWR VGND sg13g2_fill_2
XFILLER_31_84 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2853_ heichips25_sap3/net70 heichips25_sap3/_0476_ heichips25_sap3/_0495_
+ heichips25_sap3/_0496_ VPWR VGND sg13g2_nor3_1
Xheichips25_sap3_fanout71 heichips25_sap3/_1746_ heichips25_sap3/net71 VPWR VGND sg13g2_buf_1
Xheichips25_sap3_fanout60 heichips25_sap3/_0830_ heichips25_sap3/net60 VPWR VGND sg13g2_buf_1
Xoutput40 net40 uo_out[5] VPWR VGND sg13g2_buf_1
Xheichips25_sap3__2784_ VGND VPWR heichips25_sap3/_1646_ heichips25_sap3/_0428_ heichips25_sap3/_0429_
+ heichips25_sap3/net221 sg13g2_a21oi_1
Xheichips25_sap3_fanout82 heichips25_sap3/_1740_ heichips25_sap3/net82 VPWR VGND sg13g2_buf_1
Xheichips25_sap3_fanout93 heichips25_sap3/_1187_ heichips25_sap3/net93 VPWR VGND sg13g2_buf_1
XFILLER_49_744 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3405_ heichips25_sap3/_1010_ heichips25_sap3/_1011_ heichips25_sap3/_1009_
+ heichips25_sap3/_1012_ VPWR VGND sg13g2_nand3_1
Xheichips25_can_lehmann_fsm__2989__669 VPWR VGND net668 sg13g2_tiehi
XFILLER_0_283 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3336_ heichips25_sap3/_0946_ heichips25_sap3/_0926_ heichips25_sap3/_0943_
+ VPWR VGND sg13g2_xnor2_1
Xheichips25_sap3__3267_ heichips25_sap3/_0314_ VPWR heichips25_sap3/_0880_ VGND heichips25_sap3/_1719_
+ heichips25_sap3/_0879_ sg13g2_o21ai_1
XFILLER_44_471 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2218_ heichips25_sap3/_1562_ heichips25_sap3/_1611_ heichips25_sap3/_1634_
+ heichips25_sap3/_1638_ heichips25_sap3/_1639_ VPWR VGND sg13g2_nor4_1
Xheichips25_sap3__3198_ heichips25_sap3/_0811_ heichips25_sap3__4006_/Q heichips25_sap3/net148
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__2149_ heichips25_sap3/_1496_ heichips25_sap3/_1568_ heichips25_sap3/_1570_
+ VPWR VGND sg13g2_nor2_1
XFILLER_9_840 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__3040_ net758 VGND VPWR heichips25_can_lehmann_fsm/net945
+ heichips25_can_lehmann_fsm__3040_/Q clknet_leaf_22_clk sg13g2_dfrbpq_1
Xclkbuf_4_9_0_heichips25_sap3\_sap_3_inst.alu_inst.clk clknet_0_heichips25_sap3\/sap_3_inst.alu_inst.clk
+ clknet_4_9_0_heichips25_sap3\/sap_3_inst.alu_inst.clk VPWR VGND sg13g2_buf_8
Xheichips25_can_lehmann_fsm__2824_ net558 VGND VPWR heichips25_can_lehmann_fsm/_0049_
+ heichips25_can_lehmann_fsm__2824_/Q clknet_leaf_10_clk sg13g2_dfrbpq_1
Xclkbuf_leaf_19_clk clknet_2_2__leaf_clk clknet_leaf_19_clk VPWR VGND sg13g2_buf_8
XFILLER_27_438 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2755_ VGND VPWR heichips25_can_lehmann_fsm/_0856_ heichips25_can_lehmann_fsm/net426
+ heichips25_can_lehmann_fsm/_0277_ heichips25_can_lehmann_fsm/_0843_ sg13g2_a21oi_1
XFILLER_36_994 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1706_ heichips25_can_lehmann_fsm/_1016_ heichips25_can_lehmann_fsm/_1029_
+ heichips25_can_lehmann_fsm/_1030_ VPWR VGND sg13g2_nor2_1
Xheichips25_can_lehmann_fsm__2686_ heichips25_can_lehmann_fsm/net468 VPWR heichips25_can_lehmann_fsm/_0809_
+ VGND heichips25_can_lehmann_fsm/net1033 heichips25_can_lehmann_fsm/net398 sg13g2_o21ai_1
XFILLER_23_655 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1637_ VPWR heichips25_can_lehmann_fsm/_0961_ heichips25_can_lehmann_fsm/net939
+ VGND sg13g2_inv_1
XFILLER_10_305 VPWR VGND sg13g2_fill_1
XFILLER_10_316 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1568_ VPWR heichips25_can_lehmann_fsm/_0892_ heichips25_can_lehmann_fsm/net978
+ VGND sg13g2_inv_1
XFILLER_10_327 VPWR VGND sg13g2_fill_2
XFILLER_10_349 VPWR VGND sg13g2_decap_8
XFILLER_2_526 VPWR VGND sg13g2_fill_2
XFILLER_45_257 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3121_ VPWR VGND heichips25_sap3/net266 heichips25_sap3/_0724_ heichips25_sap3/_0654_
+ heichips25_sap3/_1513_ heichips25_sap3/_0734_ heichips25_sap3/_0638_ sg13g2_a221oi_1
XFILLER_14_611 VPWR VGND sg13g2_decap_4
XFILLER_42_975 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3052_ VGND VPWR heichips25_sap3/net241 heichips25_sap3/_0659_ heichips25_sap3/_0665_
+ heichips25_sap3/_0663_ sg13g2_a21oi_1
XFILLER_26_95 VPWR VGND sg13g2_decap_8
XFILLER_42_986 VPWR VGND sg13g2_fill_2
XFILLER_9_147 VPWR VGND sg13g2_decap_8
Xclkbuf_5_18__f_heichips25_sap3\_sap_3_inst.alu_inst.clk heichips25_sap3__3927_/CLK
+ clknet_4_9_0_heichips25_sap3\/sap_3_inst.alu_inst.clk VPWR VGND sg13g2_buf_16
XFILLER_10_861 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3954_ heichips25_sap3/net440 VGND VPWR heichips25_sap3/_0095_ heichips25_sap3__3954_/Q
+ heichips25_sap3__4016_/CLK sg13g2_dfrbpq_1
Xheichips25_sap3__3885_ heichips25_sap3/net451 VGND VPWR heichips25_sap3/_0026_ heichips25_sap3__3885_/Q
+ heichips25_sap3__3921_/CLK sg13g2_dfrbpq_1
XFILLER_5_353 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__2905_ heichips25_sap3/_0380_ heichips25_sap3/_0368_ heichips25_sap3/_0545_
+ VPWR VGND sg13g2_xor2_1
Xheichips25_sap3__2836_ heichips25_sap3/_0478_ VPWR heichips25_sap3/_0479_ VGND heichips25_sap3/net284
+ heichips25_sap3/_0441_ sg13g2_o21ai_1
XFILLER_3_11 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2767_ heichips25_sap3/_0399_ heichips25_sap3/_0409_ heichips25_sap3/_0412_
+ heichips25_sap3/_0413_ VPWR VGND sg13g2_nor3_1
Xheichips25_sap3__2698_ heichips25_sap3/_1896_ heichips25_sap3/_0213_ heichips25_sap3/_0342_
+ heichips25_sap3/net154 heichips25_sap3/_0344_ VPWR VGND sg13g2_nor4_1
XFILLER_3_88 VPWR VGND sg13g2_decap_8
XFILLER_3_77 VPWR VGND sg13g2_decap_4
XFILLER_3_1028 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3319_ heichips25_sap3/_0930_ heichips25_sap3/net68 uio_oe_sap3\[2\]
+ VPWR VGND sg13g2_nand2b_1
Xheichips25_can_lehmann_fsm__2540_ heichips25_can_lehmann_fsm/net466 VPWR heichips25_can_lehmann_fsm/_0736_
+ VGND heichips25_can_lehmann_fsm/net969 heichips25_can_lehmann_fsm/net356 sg13g2_o21ai_1
XFILLER_18_983 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2471_ VGND VPWR heichips25_can_lehmann_fsm/_0930_ heichips25_can_lehmann_fsm/net418
+ heichips25_can_lehmann_fsm/_0135_ heichips25_can_lehmann_fsm/_0701_ sg13g2_a21oi_1
Xclkbuf_leaf_8_clk clknet_2_3__leaf_clk clknet_leaf_8_clk VPWR VGND sg13g2_buf_8
XFILLER_8_191 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__3023_ net698 VGND VPWR heichips25_can_lehmann_fsm/net850
+ heichips25_can_lehmann_fsm__3023_/Q clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_41_1001 VPWR VGND sg13g2_fill_2
XFILLER_27_235 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2807_ net592 VGND VPWR heichips25_can_lehmann_fsm/net1211
+ heichips25_can_lehmann_fsm__2807_/Q clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_28_769 VPWR VGND sg13g2_fill_1
XFILLER_43_728 VPWR VGND sg13g2_fill_2
XFILLER_36_791 VPWR VGND sg13g2_fill_2
XFILLER_42_238 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2738_ heichips25_can_lehmann_fsm/net470 VPWR heichips25_can_lehmann_fsm/_0835_
+ VGND heichips25_can_lehmann_fsm/net343 heichips25_can_lehmann_fsm/net355 sg13g2_o21ai_1
XFILLER_24_964 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2669_ VGND VPWR heichips25_can_lehmann_fsm/_0878_ heichips25_can_lehmann_fsm/net375
+ heichips25_can_lehmann_fsm/_0234_ heichips25_can_lehmann_fsm/_0800_ sg13g2_a21oi_1
XFILLER_11_614 VPWR VGND sg13g2_fill_1
XFILLER_24_997 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_hold868 heichips25_can_lehmann_fsm__3009_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net867 sg13g2_dlygate4sd3_1
XFILLER_10_124 VPWR VGND sg13g2_decap_8
XFILLER_11_647 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm_hold857 heichips25_can_lehmann_fsm/_0223_ VPWR VGND heichips25_can_lehmann_fsm/net856
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold846 heichips25_can_lehmann_fsm/_0225_ VPWR VGND heichips25_can_lehmann_fsm/net845
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold879 heichips25_can_lehmann_fsm/_0268_ VPWR VGND heichips25_can_lehmann_fsm/net878
+ sg13g2_dlygate4sd3_1
XFILLER_6_139 VPWR VGND sg13g2_decap_8
XFILLER_10_179 VPWR VGND sg13g2_decap_4
XFILLER_12_53 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3670_ heichips25_sap3/_0888_ VPWR heichips25_sap3/_1214_ VGND heichips25_sap3/net111
+ heichips25_sap3/_1213_ sg13g2_o21ai_1
Xheichips25_sap3__2621_ heichips25_sap3/_1360_ heichips25_sap3/net835 heichips25_sap3/_0290_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_can_lehmann_fsm__2951__532 VPWR VGND net531 sg13g2_tiehi
XFILLER_2_389 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2552_ heichips25_sap3/_0225_ heichips25_sap3/_0226_ heichips25_sap3/_0227_
+ VPWR VGND sg13g2_and2_1
Xheichips25_sap3__2483_ heichips25_sap3/_1880_ heichips25_sap3/_1882_ heichips25_sap3/_1896_
+ VPWR VGND sg13g2_nor2_1
XFILLER_46_533 VPWR VGND sg13g2_fill_1
XFILLER_37_94 VPWR VGND sg13g2_fill_1
XFILLER_37_83 VPWR VGND sg13g2_fill_1
XFILLER_18_235 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3104_ heichips25_sap3/_0717_ heichips25_sap3/_0714_ heichips25_sap3/_0716_
+ VPWR VGND sg13g2_nand2_1
XFILLER_26_290 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3035_ VGND VPWR heichips25_sap3/_1486_ heichips25_sap3/_1572_ heichips25_sap3/_0648_
+ heichips25_sap3/_1510_ sg13g2_a21oi_1
XFILLER_41_271 VPWR VGND sg13g2_decap_8
XFILLER_14_485 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3937_ heichips25_sap3/net441 VGND VPWR heichips25_sap3/_0078_ heichips25_sap3__3937_/Q
+ clkload20/A sg13g2_dfrbpq_1
Xheichips25_sap3__3868_ heichips25_sap3__3887_/Q heichips25_sap3/net1124 heichips25_sap3/_0007_
+ heichips25_sap3/_0195_ VPWR VGND sg13g2_mux2_1
Xheichips25_sap3__2819_ heichips25_sap3/_1870_ VPWR heichips25_sap3/_0463_ VGND heichips25_sap3/net288
+ heichips25_sap3/_0462_ sg13g2_o21ai_1
Xheichips25_sap3__3799_ heichips25_sap3/_1305_ heichips25_sap3/_1306_ heichips25_sap3/_1304_
+ heichips25_sap3/_1308_ VPWR VGND heichips25_sap3/_1307_ sg13g2_nand4_1
Xheichips25_can_lehmann_fsm__2930__616 VPWR VGND net615 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__1971_ VGND VPWR heichips25_can_lehmann_fsm/net345 heichips25_can_lehmann_fsm/net192
+ heichips25_can_lehmann_fsm/_0331_ heichips25_can_lehmann_fsm/net181 sg13g2_a21oi_1
XFILLER_49_382 VPWR VGND sg13g2_decap_4
XFILLER_25_739 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2523_ VGND VPWR heichips25_can_lehmann_fsm/_0917_ heichips25_can_lehmann_fsm/net415
+ heichips25_can_lehmann_fsm/_0161_ heichips25_can_lehmann_fsm/_0727_ sg13g2_a21oi_1
XFILLER_33_761 VPWR VGND sg13g2_decap_8
XFILLER_21_956 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2454_ heichips25_can_lehmann_fsm/net472 VPWR heichips25_can_lehmann_fsm/_0693_
+ VGND heichips25_can_lehmann_fsm/net1024 heichips25_can_lehmann_fsm/net404 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2385_ VGND VPWR heichips25_can_lehmann_fsm/_0955_ heichips25_can_lehmann_fsm/net372
+ heichips25_can_lehmann_fsm/_0092_ heichips25_can_lehmann_fsm/_0658_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__3006_ net545 VGND VPWR heichips25_can_lehmann_fsm/net932
+ heichips25_can_lehmann_fsm__3006_/Q clknet_leaf_15_clk sg13g2_dfrbpq_1
XFILLER_0_838 VPWR VGND sg13g2_fill_2
XFILLER_28_566 VPWR VGND sg13g2_fill_2
XFILLER_23_260 VPWR VGND sg13g2_fill_1
XFILLER_7_404 VPWR VGND sg13g2_decap_4
XFILLER_48_1007 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__1983_ VPWR heichips25_sap3/_1409_ heichips25_sap3__3968_/Q VGND
+ sg13g2_inv_1
Xheichips25_sap3__3722_ heichips25_sap3__4023_/Q heichips25_sap3/_1138_ heichips25_sap3/net117
+ heichips25_sap3/_0164_ VPWR VGND sg13g2_mux2_1
XFILLER_3_621 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3653_ heichips25_sap3/_1201_ heichips25_sap3/_0327_ heichips25_sap3/net146
+ heichips25_sap3/_1200_ VPWR VGND sg13g2_and3_1
Xheichips25_sap3__2604_ heichips25_sap3/_0276_ heichips25_sap3/_0272_ heichips25_sap3/_0275_
+ VPWR VGND sg13g2_xnor2_1
Xheichips25_sap3__3584_ heichips25_sap3/_1161_ heichips25_sap3/net95 net46 VPWR VGND
+ sg13g2_nand2b_1
Xheichips25_sap3__2535_ heichips25_sap3/_0199_ heichips25_sap3/_0200_ heichips25_sap3/_0203_
+ heichips25_sap3/_0211_ uio_out_sap3\[0\] VPWR VGND sg13g2_or4_1
Xheichips25_sap3__2466_ heichips25_sap3/_1865_ VPWR heichips25_sap3/_1879_ VGND heichips25_sap3/net224
+ heichips25_sap3/_1874_ sg13g2_o21ai_1
XFILLER_47_897 VPWR VGND sg13g2_fill_1
XFILLER_34_514 VPWR VGND sg13g2_decap_8
XFILLER_19_599 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__2397_ heichips25_sap3/_1815_ VPWR heichips25_sap3/_1816_ VGND heichips25_sap3/net277
+ heichips25_sap3/net155 sg13g2_o21ai_1
XFILLER_21_208 VPWR VGND sg13g2_decap_8
XFILLER_15_794 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2860__776 VPWR VGND net775 sg13g2_tiehi
XFILLER_9_76 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3018_ heichips25_sap3/net232 uio_out_sap3\[4\] heichips25_sap3/_0635_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_can_lehmann_fsm__2170_ heichips25_can_lehmann_fsm/_0507_ heichips25_can_lehmann_fsm/_0506_
+ heichips25_can_lehmann_fsm/_1097_ VPWR VGND sg13g2_nand2b_1
XFILLER_6_470 VPWR VGND sg13g2_decap_8
Xclkbuf_5_1__f_heichips25_sap3\_sap_3_inst.alu_inst.clk heichips25_sap3__3996_/CLK
+ clknet_4_0_0_heichips25_sap3\/sap_3_inst.alu_inst.clk VPWR VGND sg13g2_buf_16
XFILLER_49_190 VPWR VGND sg13g2_fill_2
XFILLER_38_864 VPWR VGND sg13g2_fill_2
XFILLER_37_330 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1954_ heichips25_can_lehmann_fsm/_1062_ heichips25_can_lehmann_fsm/net1253
+ heichips25_can_lehmann_fsm/_0316_ VPWR VGND sg13g2_xor2_1
XFILLER_37_363 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1885_ heichips25_can_lehmann_fsm/_1176_ heichips25_can_lehmann_fsm/_1198_
+ heichips25_can_lehmann_fsm/_0002_ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3_fanout436 heichips25_sap3/net437 heichips25_sap3/net436 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout447 heichips25_sap3/net449 heichips25_sap3/net447 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout458 heichips25_sap3/net462 heichips25_sap3/net458 VPWR VGND
+ sg13g2_buf_1
XFILLER_40_539 VPWR VGND sg13g2_fill_2
XFILLER_33_591 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2906__684 VPWR VGND net683 sg13g2_tiehi
Xheichips25_can_lehmann_fsm__2506_ heichips25_can_lehmann_fsm/net491 VPWR heichips25_can_lehmann_fsm/_0719_
+ VGND heichips25_can_lehmann_fsm__2928_/Q heichips25_can_lehmann_fsm/net421 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm__2437_ VGND VPWR heichips25_can_lehmann_fsm/_0938_ heichips25_can_lehmann_fsm/net368
+ heichips25_can_lehmann_fsm/_0118_ heichips25_can_lehmann_fsm/_0684_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__2368_ heichips25_can_lehmann_fsm/net501 VPWR heichips25_can_lehmann_fsm/_0650_
+ VGND heichips25_can_lehmann_fsm__2858_/Q heichips25_can_lehmann_fsm/net387 sg13g2_o21ai_1
XFILLER_20_285 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2299_ heichips25_can_lehmann_fsm/net327 VPWR heichips25_can_lehmann_fsm/_0610_
+ VGND heichips25_can_lehmann_fsm/net983 heichips25_can_lehmann_fsm/_0607_ sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm_fanout373 heichips25_can_lehmann_fsm/net389 heichips25_can_lehmann_fsm/net373
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout362 heichips25_can_lehmann_fsm/net389 heichips25_can_lehmann_fsm/net362
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout351 heichips25_can_lehmann_fsm__2776_/Q heichips25_can_lehmann_fsm/net351
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout384 heichips25_can_lehmann_fsm/net387 heichips25_can_lehmann_fsm/net384
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout395 heichips25_can_lehmann_fsm/net397 heichips25_can_lehmann_fsm/net395
+ VPWR VGND sg13g2_buf_1
Xheichips25_sap3__2320_ heichips25_sap3/_1694_ heichips25_sap3/_1713_ heichips25_sap3/_1732_
+ heichips25_sap3/_1741_ VPWR VGND sg13g2_nor3_1
Xheichips25_sap3__2251_ heichips25_sap3/_1574_ heichips25_sap3/_1670_ heichips25_sap3/_1671_
+ heichips25_sap3/_1672_ VPWR VGND sg13g2_nor3_1
XFILLER_28_374 VPWR VGND sg13g2_decap_4
XFILLER_29_897 VPWR VGND sg13g2_fill_1
XFILLER_43_333 VPWR VGND sg13g2_fill_2
XFILLER_43_322 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2182_ heichips25_sap3/_1548_ heichips25_sap3/_1602_ heichips25_sap3/net229
+ heichips25_sap3/_1603_ VPWR VGND sg13g2_nand3_1
XFILLER_11_241 VPWR VGND sg13g2_fill_2
XFILLER_15_1017 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__2807__593 VPWR VGND net592 sg13g2_tiehi
Xheichips25_sap3__1966_ VPWR heichips25_sap3/_1392_ heichips25_sap3__3931_/Q VGND
+ sg13g2_inv_1
XFILLER_3_440 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3705_ heichips25_sap3/_0154_ heichips25_sap3/_0929_ heichips25_sap3/_1235_
+ heichips25_sap3/net115 heichips25_sap3/_1376_ VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__3636_ heichips25_sap3/_1066_ heichips25_sap3__3989_/Q heichips25_sap3/net93
+ heichips25_sap3/_0130_ VPWR VGND sg13g2_mux2_1
Xheichips25_sap3__3874__819 VPWR net818 heichips25_sap3__4021_/CLK VGND sg13g2_inv_1
Xheichips25_sap3__3567_ heichips25_sap3/_1055_ heichips25_sap3/_1086_ heichips25_sap3/_1146_
+ heichips25_sap3/_1147_ heichips25_sap3/_1148_ VPWR VGND sg13g2_nor4_1
Xheichips25_sap3__3498_ heichips25_sap3/net119 heichips25_sap3/_0901_ heichips25_sap3/_1094_
+ VPWR VGND sg13g2_nor2_1
Xheichips25_sap3__2518_ heichips25_sap3/_1929_ heichips25_sap3/net76 heichips25_sap3__3979_/Q
+ heichips25_sap3/net83 heichips25_sap3__3955_/Q VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3__2449_ heichips25_sap3/_1863_ heichips25_sap3/_1859_ heichips25_sap3/net66
+ heichips25_sap3/_1864_ VPWR VGND sg13g2_a21o_1
XFILLER_34_300 VPWR VGND sg13g2_fill_2
XFILLER_46_171 VPWR VGND sg13g2_decap_4
XFILLER_35_867 VPWR VGND sg13g2_fill_1
XFILLER_35_834 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1670_ heichips25_can_lehmann_fsm/net350 heichips25_can_lehmann_fsm/_0992_
+ heichips25_can_lehmann_fsm/_0994_ VPWR VGND sg13g2_and2_1
XFILLER_22_517 VPWR VGND sg13g2_fill_2
XFILLER_30_583 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2222_ heichips25_can_lehmann_fsm/_0548_ heichips25_can_lehmann_fsm/_0547_
+ heichips25_can_lehmann_fsm/_1105_ VPWR VGND sg13g2_nand2b_1
Xheichips25_can_lehmann_fsm__2153_ heichips25_can_lehmann_fsm/_0491_ heichips25_can_lehmann_fsm/_0490_
+ heichips25_can_lehmann_fsm/_0489_ heichips25_can_lehmann_fsm/_0492_ VPWR VGND sg13g2_a21o_1
Xheichips25_can_lehmann_fsm__2084_ heichips25_can_lehmann_fsm/_0427_ heichips25_can_lehmann_fsm/net345
+ heichips25_can_lehmann_fsm/_1056_ VPWR VGND sg13g2_xnor2_1
Xheichips25_can_lehmann_fsm__2986_ net680 VGND VPWR heichips25_can_lehmann_fsm/net979
+ heichips25_can_lehmann_fsm__2986_/Q clknet_leaf_18_clk sg13g2_dfrbpq_1
XFILLER_44_108 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm__1937_ VGND VPWR heichips25_can_lehmann_fsm__2954_/Q heichips25_can_lehmann_fsm/net308
+ heichips25_can_lehmann_fsm/_0300_ heichips25_can_lehmann_fsm/_0299_ sg13g2_a21oi_1
Xheichips25_sap3_fanout211 heichips25_sap3/net212 heichips25_sap3/net211 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout222 heichips25_sap3/_1625_ heichips25_sap3/net222 VPWR VGND
+ sg13g2_buf_1
XFILLER_25_333 VPWR VGND sg13g2_fill_2
XFILLER_26_834 VPWR VGND sg13g2_decap_8
Xheichips25_sap3_fanout244 heichips25_sap3/_1512_ heichips25_sap3/net244 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout255 heichips25_sap3/_1488_ heichips25_sap3/net255 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout266 heichips25_sap3__3926_/Q heichips25_sap3/net266 VPWR VGND
+ sg13g2_buf_1
Xheichips25_can_lehmann_fsm__1868_ heichips25_can_lehmann_fsm/_1182_ VPWR heichips25_can_lehmann_fsm/_1183_
+ VGND heichips25_can_lehmann_fsm__2867_/Q heichips25_can_lehmann_fsm/net335 sg13g2_o21ai_1
Xheichips25_sap3_fanout233 heichips25_sap3/_1466_ heichips25_sap3/net233 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout288 heichips25_sap3/net289 heichips25_sap3/net288 VPWR VGND
+ sg13g2_buf_1
Xheichips25_sap3_fanout277 heichips25_sap3__3905_/Q heichips25_sap3/net277 VPWR VGND
+ sg13g2_buf_1
Xheichips25_can_lehmann_fsm__2982__697 VPWR VGND net696 sg13g2_tiehi
XFILLER_25_399 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm__1799_ heichips25_can_lehmann_fsm/_0886_ heichips25_can_lehmann_fsm/_0991_
+ heichips25_can_lehmann_fsm/_1115_ VPWR VGND sg13g2_nor2_1
XFILLER_40_336 VPWR VGND sg13g2_decap_8
XFILLER_5_716 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm_fanout170 heichips25_can_lehmann_fsm/net174 heichips25_can_lehmann_fsm/net170
+ VPWR VGND sg13g2_buf_1
Xheichips25_can_lehmann_fsm_fanout181 heichips25_can_lehmann_fsm/_0312_ heichips25_can_lehmann_fsm/net181
+ VPWR VGND sg13g2_buf_1
XFILLER_1_933 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm_fanout192 heichips25_can_lehmann_fsm/net194 heichips25_can_lehmann_fsm/net192
+ VPWR VGND sg13g2_buf_1
Xheichips25_sap3__3421_ net43 uio_oe_sap3\[6\] heichips25_sap3/net68 heichips25_sap3/_1028_
+ VPWR VGND sg13g2_mux2_1
XFILLER_0_498 VPWR VGND sg13g2_decap_8
Xheichips25_sap3__3352_ heichips25_sap3/_0961_ heichips25_sap3/net132 heichips25_sap3__3991_/Q
+ heichips25_sap3/net142 heichips25_sap3__3983_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_35_108 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2303_ heichips25_sap3/_1536_ heichips25_sap3/_1572_ heichips25_sap3/_1724_
+ VPWR VGND sg13g2_nor2_1
XFILLER_21_1021 VPWR VGND sg13g2_decap_8
XFILLER_17_845 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3283_ VPWR VGND heichips25_sap3__3940_/Q heichips25_sap3/_0894_
+ heichips25_sap3/net105 heichips25_sap3__3948_/Q heichips25_sap3/_0895_ heichips25_sap3/net108
+ sg13g2_a221oi_1
Xheichips25_sap3__2234_ heichips25_sap3/_1655_ heichips25_sap3/net268 heichips25_sap3/_1501_
+ VPWR VGND sg13g2_nand2_1
XFILLER_43_185 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__2165_ heichips25_sap3/_1574_ heichips25_sap3/_1583_ heichips25_sap3/_1586_
+ VPWR VGND sg13g2_nor2_1
XFILLER_32_826 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2096_ heichips25_sap3/_1506_ heichips25_sap3/_1511_ heichips25_sap3/_1517_
+ VPWR VGND sg13g2_nor2_1
XFILLER_6_55 VPWR VGND sg13g2_decap_4
XFILLER_4_760 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2998_ heichips25_sap3/_0626_ uio_out_sap3\[1\] heichips25_sap3/net201
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__1949_ VPWR heichips25_sap3/_1375_ heichips25_sap3__3933_/Q VGND
+ sg13g2_inv_1
Xheichips25_sap3__3619_ heichips25_sap3/_0122_ heichips25_sap3/_0929_ heichips25_sap3/_1181_
+ heichips25_sap3/net102 heichips25_sap3/_1378_ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2840_ net526 VGND VPWR heichips25_can_lehmann_fsm/_0065_
+ heichips25_can_lehmann_fsm__2840_/Q clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_13_2 VPWR VGND sg13g2_fill_1
XFILLER_47_480 VPWR VGND sg13g2_decap_4
Xheichips25_can_lehmann_fsm__2771_ VGND VPWR heichips25_can_lehmann_fsm/_0852_ heichips25_can_lehmann_fsm/net400
+ heichips25_can_lehmann_fsm/_0285_ heichips25_can_lehmann_fsm/_0851_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm__1722_ heichips25_can_lehmann_fsm/net1195 heichips25_can_lehmann_fsm/net1174
+ heichips25_can_lehmann_fsm__2818_/Q heichips25_can_lehmann_fsm/_1043_ VPWR VGND
+ sg13g2_nor3_1
XFILLER_34_152 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1653_ VPWR heichips25_can_lehmann_fsm/_0977_ heichips25_can_lehmann_fsm/net1255
+ VGND sg13g2_inv_1
XFILLER_34_174 VPWR VGND sg13g2_decap_8
XFILLER_34_185 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__1584_ VPWR heichips25_can_lehmann_fsm/_0908_ heichips25_can_lehmann_fsm/net1103
+ VGND sg13g2_inv_1
Xheichips25_can_lehmann_fsm__2205_ heichips25_can_lehmann_fsm/_0535_ heichips25_can_lehmann_fsm/net165
+ heichips25_can_lehmann_fsm/_0534_ heichips25_can_lehmann_fsm/net175 heichips25_can_lehmann_fsm/net851
+ VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm__2136_ heichips25_can_lehmann_fsm__3048_/Q heichips25_can_lehmann_fsm/_0474_
+ heichips25_can_lehmann_fsm/_1162_ heichips25_can_lehmann_fsm/_0475_ VPWR VGND sg13g2_mux2_1
Xheichips25_can_lehmann_fsm__2067_ VPWR VGND heichips25_can_lehmann_fsm/_0413_ heichips25_can_lehmann_fsm/_1176_
+ heichips25_can_lehmann_fsm/_0412_ heichips25_can_lehmann_fsm/_0977_ heichips25_can_lehmann_fsm/_0019_
+ heichips25_can_lehmann_fsm/net181 sg13g2_a221oi_1
XFILLER_46_929 VPWR VGND sg13g2_fill_1
Xheichips25_can_lehmann_fsm__2969_ net748 VGND VPWR heichips25_can_lehmann_fsm/_0194_
+ heichips25_can_lehmann_fsm__2969_/Q clknet_leaf_20_clk sg13g2_dfrbpq_1
XFILLER_13_325 VPWR VGND sg13g2_fill_1
XFILLER_14_848 VPWR VGND sg13g2_fill_2
Xheichips25_can_lehmann_fsm_hold1175 heichips25_can_lehmann_fsm__2819_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1174 sg13g2_dlygate4sd3_1
XFILLER_15_97 VPWR VGND sg13g2_decap_8
Xheichips25_can_lehmann_fsm_hold1153 heichips25_can_lehmann_fsm__3028_/Q VPWR VGND
+ heichips25_can_lehmann_fsm/net1152 sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1197 heichips25_can_lehmann_fsm/_0045_ VPWR VGND heichips25_can_lehmann_fsm/net1196
+ sg13g2_dlygate4sd3_1
Xheichips25_can_lehmann_fsm_hold1186 heichips25_can_lehmann_fsm/_0047_ VPWR VGND heichips25_can_lehmann_fsm/net1185
+ sg13g2_dlygate4sd3_1
Xheichips25_sap3__3970_ heichips25_sap3/net440 VGND VPWR heichips25_sap3/_0111_ heichips25_sap3__3970_/Q
+ heichips25_sap3__4018_/CLK sg13g2_dfrbpq_1
Xheichips25_sap3_hold840 heichips25_sap3/_0185_ VPWR VGND heichips25_sap3/net839 sg13g2_dlygate4sd3_1
Xheichips25_sap3__2921_ net43 heichips25_sap3/net157 heichips25_sap3/_0560_ VPWR VGND
+ sg13g2_nor2b_1
XFILLER_31_41 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2852_ VPWR VGND heichips25_sap3/_0494_ heichips25_sap3/net158 heichips25_sap3/_0493_
+ heichips25_sap3__3909_/Q heichips25_sap3/_0495_ heichips25_sap3/net204 sg13g2_a221oi_1
Xheichips25_sap3_fanout72 heichips25_sap3/_1746_ heichips25_sap3/net72 VPWR VGND sg13g2_buf_1
Xheichips25_sap3_fanout50 heichips25_sap3/_0922_ heichips25_sap3/net50 VPWR VGND sg13g2_buf_1
Xheichips25_sap3_fanout61 heichips25_sap3/net62 heichips25_sap3/net61 VPWR VGND sg13g2_buf_1
Xoutput41 net41 uo_out[6] VPWR VGND sg13g2_buf_1
Xheichips25_sap3__2783_ heichips25_sap3/_1761_ heichips25_sap3/_0426_ heichips25_sap3/_1755_
+ heichips25_sap3/_0428_ VPWR VGND heichips25_sap3/_0427_ sg13g2_nand4_1
Xoutput30 net30 uio_out[3] VPWR VGND sg13g2_buf_1
Xheichips25_sap3_fanout83 heichips25_sap3/_1739_ heichips25_sap3/net83 VPWR VGND sg13g2_buf_1
Xheichips25_sap3_fanout94 heichips25_sap3/_1171_ heichips25_sap3/net94 VPWR VGND sg13g2_buf_1
XFILLER_49_734 VPWR VGND sg13g2_decap_4
XFILLER_49_723 VPWR VGND sg13g2_decap_4
Xheichips25_sap3__3404_ heichips25_sap3/_1011_ heichips25_sap3/_0768_ heichips25_sap3__3977_/Q
+ heichips25_sap3/net143 heichips25_sap3__3985_/Q VPWR VGND sg13g2_a22oi_1
XFILLER_48_299 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__3335_ VPWR heichips25_sap3/_0945_ heichips25_sap3/_0944_ VGND sg13g2_inv_1
Xheichips25_sap3__3266_ VGND VPWR heichips25_sap3/_0707_ heichips25_sap3/_0878_ heichips25_sap3/_0879_
+ heichips25_sap3/_0699_ sg13g2_a21oi_1
XFILLER_45_995 VPWR VGND sg13g2_fill_2
Xheichips25_sap3__2217_ heichips25_sap3/_1638_ heichips25_sap3/_1637_ heichips25_sap3/_1571_
+ VPWR VGND sg13g2_nand2b_1
Xheichips25_can_lehmann_fsm__2926__632 VPWR VGND net631 sg13g2_tiehi
XFILLER_44_494 VPWR VGND sg13g2_fill_1
Xheichips25_sap3__3197_ heichips25_sap3/_0808_ heichips25_sap3/_0809_ heichips25_sap3/_0807_
+ heichips25_sap3/_0810_ VPWR VGND sg13g2_nand3_1
Xheichips25_sap3__2148_ heichips25_sap3/_1569_ heichips25_sap3/_1546_ heichips25_sap3/_1566_
+ VPWR VGND sg13g2_nand2_1
Xheichips25_sap3__2079_ heichips25_sap3/_1493_ VPWR heichips25_sap3/_1500_ VGND heichips25_sap3/_1495_
+ heichips25_sap3/_1498_ sg13g2_o21ai_1
XFILLER_8_351 VPWR VGND sg13g2_decap_8
.ends

