module heichips25_tiny_wrapper2 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00_;
 wire _01_;
 wire clknet_leaf_1_clk;
 wire net525;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire \uio_oe_sap3[0] ;
 wire \uio_oe_sap3[1] ;
 wire \uio_oe_sap3[2] ;
 wire \uio_oe_sap3[3] ;
 wire \uio_oe_sap3[4] ;
 wire \uio_oe_sap3[5] ;
 wire \uio_oe_sap3[6] ;
 wire \uio_oe_sap3[7] ;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire \uio_out_sap3[0] ;
 wire \uio_out_sap3[1] ;
 wire \uio_out_sap3[2] ;
 wire \uio_out_sap3[3] ;
 wire \uio_out_sap3[4] ;
 wire \uio_out_sap3[5] ;
 wire \uio_out_sap3[6] ;
 wire \uio_out_sap3[7] ;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire \uo_out_fsm[0] ;
 wire \uo_out_fsm[1] ;
 wire \uo_out_fsm[2] ;
 wire \uo_out_fsm[3] ;
 wire \uo_out_fsm[4] ;
 wire \uo_out_fsm[5] ;
 wire \uo_out_fsm[6] ;
 wire \uo_out_fsm[7] ;
 wire \uo_out_sap3[0] ;
 wire \uo_out_sap3[1] ;
 wire \uo_out_sap3[2] ;
 wire \uo_out_sap3[3] ;
 wire \uo_out_sap3[4] ;
 wire \uo_out_sap3[5] ;
 wire net524;
 wire clknet_leaf_2_clk;
 wire \heichips25_can_lehmann_fsm/_0000_ ;
 wire \heichips25_can_lehmann_fsm/_0001_ ;
 wire \heichips25_can_lehmann_fsm/_0002_ ;
 wire \heichips25_can_lehmann_fsm/_0003_ ;
 wire \heichips25_can_lehmann_fsm/_0004_ ;
 wire \heichips25_can_lehmann_fsm/_0005_ ;
 wire \heichips25_can_lehmann_fsm/_0006_ ;
 wire \heichips25_can_lehmann_fsm/_0007_ ;
 wire \heichips25_can_lehmann_fsm/_0008_ ;
 wire \heichips25_can_lehmann_fsm/_0009_ ;
 wire \heichips25_can_lehmann_fsm/_0010_ ;
 wire \heichips25_can_lehmann_fsm/_0011_ ;
 wire \heichips25_can_lehmann_fsm/_0012_ ;
 wire \heichips25_can_lehmann_fsm/_0013_ ;
 wire \heichips25_can_lehmann_fsm/_0014_ ;
 wire \heichips25_can_lehmann_fsm/_0015_ ;
 wire \heichips25_can_lehmann_fsm/_0016_ ;
 wire \heichips25_can_lehmann_fsm/_0017_ ;
 wire \heichips25_can_lehmann_fsm/_0018_ ;
 wire \heichips25_can_lehmann_fsm/_0019_ ;
 wire \heichips25_can_lehmann_fsm/_0020_ ;
 wire \heichips25_can_lehmann_fsm/_0021_ ;
 wire \heichips25_can_lehmann_fsm/_0022_ ;
 wire \heichips25_can_lehmann_fsm/_0023_ ;
 wire \heichips25_can_lehmann_fsm/_0024_ ;
 wire \heichips25_can_lehmann_fsm/_0025_ ;
 wire \heichips25_can_lehmann_fsm/_0026_ ;
 wire \heichips25_can_lehmann_fsm/_0027_ ;
 wire \heichips25_can_lehmann_fsm/_0028_ ;
 wire \heichips25_can_lehmann_fsm/_0029_ ;
 wire \heichips25_can_lehmann_fsm/_0030_ ;
 wire \heichips25_can_lehmann_fsm/_0031_ ;
 wire \heichips25_can_lehmann_fsm/_0032_ ;
 wire \heichips25_can_lehmann_fsm/_0033_ ;
 wire \heichips25_can_lehmann_fsm/_0034_ ;
 wire \heichips25_can_lehmann_fsm/_0035_ ;
 wire \heichips25_can_lehmann_fsm/_0036_ ;
 wire \heichips25_can_lehmann_fsm/_0037_ ;
 wire \heichips25_can_lehmann_fsm/_0038_ ;
 wire \heichips25_can_lehmann_fsm/_0039_ ;
 wire \heichips25_can_lehmann_fsm/_0040_ ;
 wire \heichips25_can_lehmann_fsm/_0041_ ;
 wire \heichips25_can_lehmann_fsm/_0042_ ;
 wire \heichips25_can_lehmann_fsm/_0043_ ;
 wire \heichips25_can_lehmann_fsm/_0044_ ;
 wire \heichips25_can_lehmann_fsm/_0045_ ;
 wire \heichips25_can_lehmann_fsm/_0046_ ;
 wire \heichips25_can_lehmann_fsm/_0047_ ;
 wire \heichips25_can_lehmann_fsm/_0048_ ;
 wire \heichips25_can_lehmann_fsm/_0049_ ;
 wire \heichips25_can_lehmann_fsm/_0050_ ;
 wire \heichips25_can_lehmann_fsm/_0051_ ;
 wire \heichips25_can_lehmann_fsm/_0052_ ;
 wire \heichips25_can_lehmann_fsm/_0053_ ;
 wire \heichips25_can_lehmann_fsm/_0054_ ;
 wire \heichips25_can_lehmann_fsm/_0055_ ;
 wire \heichips25_can_lehmann_fsm/_0056_ ;
 wire \heichips25_can_lehmann_fsm/_0057_ ;
 wire \heichips25_can_lehmann_fsm/_0058_ ;
 wire \heichips25_can_lehmann_fsm/_0059_ ;
 wire \heichips25_can_lehmann_fsm/_0060_ ;
 wire \heichips25_can_lehmann_fsm/_0061_ ;
 wire \heichips25_can_lehmann_fsm/_0062_ ;
 wire \heichips25_can_lehmann_fsm/_0063_ ;
 wire \heichips25_can_lehmann_fsm/_0064_ ;
 wire \heichips25_can_lehmann_fsm/_0065_ ;
 wire \heichips25_can_lehmann_fsm/_0066_ ;
 wire \heichips25_can_lehmann_fsm/_0067_ ;
 wire \heichips25_can_lehmann_fsm/_0068_ ;
 wire \heichips25_can_lehmann_fsm/_0069_ ;
 wire \heichips25_can_lehmann_fsm/_0070_ ;
 wire \heichips25_can_lehmann_fsm/_0071_ ;
 wire \heichips25_can_lehmann_fsm/_0072_ ;
 wire \heichips25_can_lehmann_fsm/_0073_ ;
 wire \heichips25_can_lehmann_fsm/_0074_ ;
 wire \heichips25_can_lehmann_fsm/_0075_ ;
 wire \heichips25_can_lehmann_fsm/_0076_ ;
 wire \heichips25_can_lehmann_fsm/_0077_ ;
 wire \heichips25_can_lehmann_fsm/_0078_ ;
 wire \heichips25_can_lehmann_fsm/_0079_ ;
 wire \heichips25_can_lehmann_fsm/_0080_ ;
 wire \heichips25_can_lehmann_fsm/_0081_ ;
 wire \heichips25_can_lehmann_fsm/_0082_ ;
 wire \heichips25_can_lehmann_fsm/_0083_ ;
 wire \heichips25_can_lehmann_fsm/_0084_ ;
 wire \heichips25_can_lehmann_fsm/_0085_ ;
 wire \heichips25_can_lehmann_fsm/_0086_ ;
 wire \heichips25_can_lehmann_fsm/_0087_ ;
 wire \heichips25_can_lehmann_fsm/_0088_ ;
 wire \heichips25_can_lehmann_fsm/_0089_ ;
 wire \heichips25_can_lehmann_fsm/_0090_ ;
 wire \heichips25_can_lehmann_fsm/_0091_ ;
 wire \heichips25_can_lehmann_fsm/_0092_ ;
 wire \heichips25_can_lehmann_fsm/_0093_ ;
 wire \heichips25_can_lehmann_fsm/_0094_ ;
 wire \heichips25_can_lehmann_fsm/_0095_ ;
 wire \heichips25_can_lehmann_fsm/_0096_ ;
 wire \heichips25_can_lehmann_fsm/_0097_ ;
 wire \heichips25_can_lehmann_fsm/_0098_ ;
 wire \heichips25_can_lehmann_fsm/_0099_ ;
 wire \heichips25_can_lehmann_fsm/_0100_ ;
 wire \heichips25_can_lehmann_fsm/_0101_ ;
 wire \heichips25_can_lehmann_fsm/_0102_ ;
 wire \heichips25_can_lehmann_fsm/_0103_ ;
 wire \heichips25_can_lehmann_fsm/_0104_ ;
 wire \heichips25_can_lehmann_fsm/_0105_ ;
 wire \heichips25_can_lehmann_fsm/_0106_ ;
 wire \heichips25_can_lehmann_fsm/_0107_ ;
 wire \heichips25_can_lehmann_fsm/_0108_ ;
 wire \heichips25_can_lehmann_fsm/_0109_ ;
 wire \heichips25_can_lehmann_fsm/_0110_ ;
 wire \heichips25_can_lehmann_fsm/_0111_ ;
 wire \heichips25_can_lehmann_fsm/_0112_ ;
 wire \heichips25_can_lehmann_fsm/_0113_ ;
 wire \heichips25_can_lehmann_fsm/_0114_ ;
 wire \heichips25_can_lehmann_fsm/_0115_ ;
 wire \heichips25_can_lehmann_fsm/_0116_ ;
 wire \heichips25_can_lehmann_fsm/_0117_ ;
 wire \heichips25_can_lehmann_fsm/_0118_ ;
 wire \heichips25_can_lehmann_fsm/_0119_ ;
 wire \heichips25_can_lehmann_fsm/_0120_ ;
 wire \heichips25_can_lehmann_fsm/_0121_ ;
 wire \heichips25_can_lehmann_fsm/_0122_ ;
 wire \heichips25_can_lehmann_fsm/_0123_ ;
 wire \heichips25_can_lehmann_fsm/_0124_ ;
 wire \heichips25_can_lehmann_fsm/_0125_ ;
 wire \heichips25_can_lehmann_fsm/_0126_ ;
 wire \heichips25_can_lehmann_fsm/_0127_ ;
 wire \heichips25_can_lehmann_fsm/_0128_ ;
 wire \heichips25_can_lehmann_fsm/_0129_ ;
 wire \heichips25_can_lehmann_fsm/_0130_ ;
 wire \heichips25_can_lehmann_fsm/_0131_ ;
 wire \heichips25_can_lehmann_fsm/_0132_ ;
 wire \heichips25_can_lehmann_fsm/_0133_ ;
 wire \heichips25_can_lehmann_fsm/_0134_ ;
 wire \heichips25_can_lehmann_fsm/_0135_ ;
 wire \heichips25_can_lehmann_fsm/_0136_ ;
 wire \heichips25_can_lehmann_fsm/_0137_ ;
 wire \heichips25_can_lehmann_fsm/_0138_ ;
 wire \heichips25_can_lehmann_fsm/_0139_ ;
 wire \heichips25_can_lehmann_fsm/_0140_ ;
 wire \heichips25_can_lehmann_fsm/_0141_ ;
 wire \heichips25_can_lehmann_fsm/_0142_ ;
 wire \heichips25_can_lehmann_fsm/_0143_ ;
 wire \heichips25_can_lehmann_fsm/_0144_ ;
 wire \heichips25_can_lehmann_fsm/_0145_ ;
 wire \heichips25_can_lehmann_fsm/_0146_ ;
 wire \heichips25_can_lehmann_fsm/_0147_ ;
 wire \heichips25_can_lehmann_fsm/_0148_ ;
 wire \heichips25_can_lehmann_fsm/_0149_ ;
 wire \heichips25_can_lehmann_fsm/_0150_ ;
 wire \heichips25_can_lehmann_fsm/_0151_ ;
 wire \heichips25_can_lehmann_fsm/_0152_ ;
 wire \heichips25_can_lehmann_fsm/_0153_ ;
 wire \heichips25_can_lehmann_fsm/_0154_ ;
 wire \heichips25_can_lehmann_fsm/_0155_ ;
 wire \heichips25_can_lehmann_fsm/_0156_ ;
 wire \heichips25_can_lehmann_fsm/_0157_ ;
 wire \heichips25_can_lehmann_fsm/_0158_ ;
 wire \heichips25_can_lehmann_fsm/_0159_ ;
 wire \heichips25_can_lehmann_fsm/_0160_ ;
 wire \heichips25_can_lehmann_fsm/_0161_ ;
 wire \heichips25_can_lehmann_fsm/_0162_ ;
 wire \heichips25_can_lehmann_fsm/_0163_ ;
 wire \heichips25_can_lehmann_fsm/_0164_ ;
 wire \heichips25_can_lehmann_fsm/_0165_ ;
 wire \heichips25_can_lehmann_fsm/_0166_ ;
 wire \heichips25_can_lehmann_fsm/_0167_ ;
 wire \heichips25_can_lehmann_fsm/_0168_ ;
 wire \heichips25_can_lehmann_fsm/_0169_ ;
 wire \heichips25_can_lehmann_fsm/_0170_ ;
 wire \heichips25_can_lehmann_fsm/_0171_ ;
 wire \heichips25_can_lehmann_fsm/_0172_ ;
 wire \heichips25_can_lehmann_fsm/_0173_ ;
 wire \heichips25_can_lehmann_fsm/_0174_ ;
 wire \heichips25_can_lehmann_fsm/_0175_ ;
 wire \heichips25_can_lehmann_fsm/_0176_ ;
 wire \heichips25_can_lehmann_fsm/_0177_ ;
 wire \heichips25_can_lehmann_fsm/_0178_ ;
 wire \heichips25_can_lehmann_fsm/_0179_ ;
 wire \heichips25_can_lehmann_fsm/_0180_ ;
 wire \heichips25_can_lehmann_fsm/_0181_ ;
 wire \heichips25_can_lehmann_fsm/_0182_ ;
 wire \heichips25_can_lehmann_fsm/_0183_ ;
 wire \heichips25_can_lehmann_fsm/_0184_ ;
 wire \heichips25_can_lehmann_fsm/_0185_ ;
 wire \heichips25_can_lehmann_fsm/_0186_ ;
 wire \heichips25_can_lehmann_fsm/_0187_ ;
 wire \heichips25_can_lehmann_fsm/_0188_ ;
 wire \heichips25_can_lehmann_fsm/_0189_ ;
 wire \heichips25_can_lehmann_fsm/_0190_ ;
 wire \heichips25_can_lehmann_fsm/_0191_ ;
 wire \heichips25_can_lehmann_fsm/_0192_ ;
 wire \heichips25_can_lehmann_fsm/_0193_ ;
 wire \heichips25_can_lehmann_fsm/_0194_ ;
 wire \heichips25_can_lehmann_fsm/_0195_ ;
 wire \heichips25_can_lehmann_fsm/_0196_ ;
 wire \heichips25_can_lehmann_fsm/_0197_ ;
 wire \heichips25_can_lehmann_fsm/_0198_ ;
 wire \heichips25_can_lehmann_fsm/_0199_ ;
 wire \heichips25_can_lehmann_fsm/_0200_ ;
 wire \heichips25_can_lehmann_fsm/_0201_ ;
 wire \heichips25_can_lehmann_fsm/_0202_ ;
 wire \heichips25_can_lehmann_fsm/_0203_ ;
 wire \heichips25_can_lehmann_fsm/_0204_ ;
 wire \heichips25_can_lehmann_fsm/_0205_ ;
 wire \heichips25_can_lehmann_fsm/_0206_ ;
 wire \heichips25_can_lehmann_fsm/_0207_ ;
 wire \heichips25_can_lehmann_fsm/_0208_ ;
 wire \heichips25_can_lehmann_fsm/_0209_ ;
 wire \heichips25_can_lehmann_fsm/_0210_ ;
 wire \heichips25_can_lehmann_fsm/_0211_ ;
 wire \heichips25_can_lehmann_fsm/_0212_ ;
 wire \heichips25_can_lehmann_fsm/_0213_ ;
 wire \heichips25_can_lehmann_fsm/_0214_ ;
 wire \heichips25_can_lehmann_fsm/_0215_ ;
 wire \heichips25_can_lehmann_fsm/_0216_ ;
 wire \heichips25_can_lehmann_fsm/_0217_ ;
 wire \heichips25_can_lehmann_fsm/_0218_ ;
 wire \heichips25_can_lehmann_fsm/_0219_ ;
 wire \heichips25_can_lehmann_fsm/_0220_ ;
 wire \heichips25_can_lehmann_fsm/_0221_ ;
 wire \heichips25_can_lehmann_fsm/_0222_ ;
 wire \heichips25_can_lehmann_fsm/_0223_ ;
 wire \heichips25_can_lehmann_fsm/_0224_ ;
 wire \heichips25_can_lehmann_fsm/_0225_ ;
 wire \heichips25_can_lehmann_fsm/_0226_ ;
 wire \heichips25_can_lehmann_fsm/_0227_ ;
 wire \heichips25_can_lehmann_fsm/_0228_ ;
 wire \heichips25_can_lehmann_fsm/_0229_ ;
 wire \heichips25_can_lehmann_fsm/_0230_ ;
 wire \heichips25_can_lehmann_fsm/_0231_ ;
 wire \heichips25_can_lehmann_fsm/_0232_ ;
 wire \heichips25_can_lehmann_fsm/_0233_ ;
 wire \heichips25_can_lehmann_fsm/_0234_ ;
 wire \heichips25_can_lehmann_fsm/_0235_ ;
 wire \heichips25_can_lehmann_fsm/_0236_ ;
 wire \heichips25_can_lehmann_fsm/_0237_ ;
 wire \heichips25_can_lehmann_fsm/_0238_ ;
 wire \heichips25_can_lehmann_fsm/_0239_ ;
 wire \heichips25_can_lehmann_fsm/_0240_ ;
 wire \heichips25_can_lehmann_fsm/_0241_ ;
 wire \heichips25_can_lehmann_fsm/_0242_ ;
 wire \heichips25_can_lehmann_fsm/_0243_ ;
 wire \heichips25_can_lehmann_fsm/_0244_ ;
 wire \heichips25_can_lehmann_fsm/_0245_ ;
 wire \heichips25_can_lehmann_fsm/_0246_ ;
 wire \heichips25_can_lehmann_fsm/_0247_ ;
 wire \heichips25_can_lehmann_fsm/_0248_ ;
 wire \heichips25_can_lehmann_fsm/_0249_ ;
 wire \heichips25_can_lehmann_fsm/_0250_ ;
 wire \heichips25_can_lehmann_fsm/_0251_ ;
 wire \heichips25_can_lehmann_fsm/_0252_ ;
 wire \heichips25_can_lehmann_fsm/_0253_ ;
 wire \heichips25_can_lehmann_fsm/_0254_ ;
 wire \heichips25_can_lehmann_fsm/_0255_ ;
 wire \heichips25_can_lehmann_fsm/_0256_ ;
 wire \heichips25_can_lehmann_fsm/_0257_ ;
 wire \heichips25_can_lehmann_fsm/_0258_ ;
 wire \heichips25_can_lehmann_fsm/_0259_ ;
 wire \heichips25_can_lehmann_fsm/_0260_ ;
 wire \heichips25_can_lehmann_fsm/_0261_ ;
 wire \heichips25_can_lehmann_fsm/_0262_ ;
 wire \heichips25_can_lehmann_fsm/_0263_ ;
 wire \heichips25_can_lehmann_fsm/_0264_ ;
 wire \heichips25_can_lehmann_fsm/_0265_ ;
 wire \heichips25_can_lehmann_fsm/_0266_ ;
 wire \heichips25_can_lehmann_fsm/_0267_ ;
 wire \heichips25_can_lehmann_fsm/_0268_ ;
 wire \heichips25_can_lehmann_fsm/_0269_ ;
 wire \heichips25_can_lehmann_fsm/_0270_ ;
 wire \heichips25_can_lehmann_fsm/_0271_ ;
 wire \heichips25_can_lehmann_fsm/_0272_ ;
 wire \heichips25_can_lehmann_fsm/_0273_ ;
 wire \heichips25_can_lehmann_fsm/_0274_ ;
 wire \heichips25_can_lehmann_fsm/_0275_ ;
 wire \heichips25_can_lehmann_fsm/_0276_ ;
 wire \heichips25_can_lehmann_fsm/_0277_ ;
 wire \heichips25_can_lehmann_fsm/_0278_ ;
 wire \heichips25_can_lehmann_fsm/_0279_ ;
 wire \heichips25_can_lehmann_fsm/_0280_ ;
 wire \heichips25_can_lehmann_fsm/_0281_ ;
 wire \heichips25_can_lehmann_fsm/_0282_ ;
 wire \heichips25_can_lehmann_fsm/_0283_ ;
 wire \heichips25_can_lehmann_fsm/_0284_ ;
 wire \heichips25_can_lehmann_fsm/_0285_ ;
 wire \heichips25_can_lehmann_fsm/_0286_ ;
 wire \heichips25_can_lehmann_fsm/_0287_ ;
 wire \heichips25_can_lehmann_fsm/_0288_ ;
 wire \heichips25_can_lehmann_fsm/_0289_ ;
 wire \heichips25_can_lehmann_fsm/_0290_ ;
 wire \heichips25_can_lehmann_fsm/_0291_ ;
 wire \heichips25_can_lehmann_fsm/_0292_ ;
 wire \heichips25_can_lehmann_fsm/_0293_ ;
 wire \heichips25_can_lehmann_fsm/_0294_ ;
 wire \heichips25_can_lehmann_fsm/_0295_ ;
 wire \heichips25_can_lehmann_fsm/_0296_ ;
 wire \heichips25_can_lehmann_fsm/_0297_ ;
 wire \heichips25_can_lehmann_fsm/_0298_ ;
 wire \heichips25_can_lehmann_fsm/_0299_ ;
 wire \heichips25_can_lehmann_fsm/_0300_ ;
 wire \heichips25_can_lehmann_fsm/_0301_ ;
 wire \heichips25_can_lehmann_fsm/_0302_ ;
 wire \heichips25_can_lehmann_fsm/_0303_ ;
 wire \heichips25_can_lehmann_fsm/_0304_ ;
 wire \heichips25_can_lehmann_fsm/_0305_ ;
 wire \heichips25_can_lehmann_fsm/_0306_ ;
 wire \heichips25_can_lehmann_fsm/_0307_ ;
 wire \heichips25_can_lehmann_fsm/_0308_ ;
 wire \heichips25_can_lehmann_fsm/_0309_ ;
 wire \heichips25_can_lehmann_fsm/_0310_ ;
 wire \heichips25_can_lehmann_fsm/_0311_ ;
 wire \heichips25_can_lehmann_fsm/_0312_ ;
 wire \heichips25_can_lehmann_fsm/_0313_ ;
 wire \heichips25_can_lehmann_fsm/_0314_ ;
 wire \heichips25_can_lehmann_fsm/_0315_ ;
 wire \heichips25_can_lehmann_fsm/_0316_ ;
 wire \heichips25_can_lehmann_fsm/_0317_ ;
 wire \heichips25_can_lehmann_fsm/_0318_ ;
 wire \heichips25_can_lehmann_fsm/_0319_ ;
 wire \heichips25_can_lehmann_fsm/_0320_ ;
 wire \heichips25_can_lehmann_fsm/_0321_ ;
 wire \heichips25_can_lehmann_fsm/_0322_ ;
 wire \heichips25_can_lehmann_fsm/_0323_ ;
 wire \heichips25_can_lehmann_fsm/_0324_ ;
 wire \heichips25_can_lehmann_fsm/_0325_ ;
 wire \heichips25_can_lehmann_fsm/_0326_ ;
 wire \heichips25_can_lehmann_fsm/_0327_ ;
 wire \heichips25_can_lehmann_fsm/_0328_ ;
 wire \heichips25_can_lehmann_fsm/_0329_ ;
 wire \heichips25_can_lehmann_fsm/_0330_ ;
 wire \heichips25_can_lehmann_fsm/_0331_ ;
 wire \heichips25_can_lehmann_fsm/_0332_ ;
 wire \heichips25_can_lehmann_fsm/_0333_ ;
 wire \heichips25_can_lehmann_fsm/_0334_ ;
 wire \heichips25_can_lehmann_fsm/_0335_ ;
 wire \heichips25_can_lehmann_fsm/_0336_ ;
 wire \heichips25_can_lehmann_fsm/_0337_ ;
 wire \heichips25_can_lehmann_fsm/_0338_ ;
 wire \heichips25_can_lehmann_fsm/_0339_ ;
 wire \heichips25_can_lehmann_fsm/_0340_ ;
 wire \heichips25_can_lehmann_fsm/_0341_ ;
 wire \heichips25_can_lehmann_fsm/_0342_ ;
 wire \heichips25_can_lehmann_fsm/_0343_ ;
 wire \heichips25_can_lehmann_fsm/_0344_ ;
 wire \heichips25_can_lehmann_fsm/_0345_ ;
 wire \heichips25_can_lehmann_fsm/_0346_ ;
 wire \heichips25_can_lehmann_fsm/_0347_ ;
 wire \heichips25_can_lehmann_fsm/_0348_ ;
 wire \heichips25_can_lehmann_fsm/_0349_ ;
 wire \heichips25_can_lehmann_fsm/_0350_ ;
 wire \heichips25_can_lehmann_fsm/_0351_ ;
 wire \heichips25_can_lehmann_fsm/_0352_ ;
 wire \heichips25_can_lehmann_fsm/_0353_ ;
 wire \heichips25_can_lehmann_fsm/_0354_ ;
 wire \heichips25_can_lehmann_fsm/_0355_ ;
 wire \heichips25_can_lehmann_fsm/_0356_ ;
 wire \heichips25_can_lehmann_fsm/_0357_ ;
 wire \heichips25_can_lehmann_fsm/_0358_ ;
 wire \heichips25_can_lehmann_fsm/_0359_ ;
 wire \heichips25_can_lehmann_fsm/_0360_ ;
 wire \heichips25_can_lehmann_fsm/_0361_ ;
 wire \heichips25_can_lehmann_fsm/_0362_ ;
 wire \heichips25_can_lehmann_fsm/_0363_ ;
 wire \heichips25_can_lehmann_fsm/_0364_ ;
 wire \heichips25_can_lehmann_fsm/_0365_ ;
 wire \heichips25_can_lehmann_fsm/_0366_ ;
 wire \heichips25_can_lehmann_fsm/_0367_ ;
 wire \heichips25_can_lehmann_fsm/_0368_ ;
 wire \heichips25_can_lehmann_fsm/_0369_ ;
 wire \heichips25_can_lehmann_fsm/_0370_ ;
 wire \heichips25_can_lehmann_fsm/_0371_ ;
 wire \heichips25_can_lehmann_fsm/_0372_ ;
 wire \heichips25_can_lehmann_fsm/_0373_ ;
 wire \heichips25_can_lehmann_fsm/_0374_ ;
 wire \heichips25_can_lehmann_fsm/_0375_ ;
 wire \heichips25_can_lehmann_fsm/_0376_ ;
 wire \heichips25_can_lehmann_fsm/_0377_ ;
 wire \heichips25_can_lehmann_fsm/_0378_ ;
 wire \heichips25_can_lehmann_fsm/_0379_ ;
 wire \heichips25_can_lehmann_fsm/_0380_ ;
 wire \heichips25_can_lehmann_fsm/_0381_ ;
 wire \heichips25_can_lehmann_fsm/_0382_ ;
 wire \heichips25_can_lehmann_fsm/_0383_ ;
 wire \heichips25_can_lehmann_fsm/_0384_ ;
 wire \heichips25_can_lehmann_fsm/_0385_ ;
 wire \heichips25_can_lehmann_fsm/_0386_ ;
 wire \heichips25_can_lehmann_fsm/_0387_ ;
 wire \heichips25_can_lehmann_fsm/_0388_ ;
 wire \heichips25_can_lehmann_fsm/_0389_ ;
 wire \heichips25_can_lehmann_fsm/_0390_ ;
 wire \heichips25_can_lehmann_fsm/_0391_ ;
 wire \heichips25_can_lehmann_fsm/_0392_ ;
 wire \heichips25_can_lehmann_fsm/_0393_ ;
 wire \heichips25_can_lehmann_fsm/_0394_ ;
 wire \heichips25_can_lehmann_fsm/_0395_ ;
 wire \heichips25_can_lehmann_fsm/_0396_ ;
 wire \heichips25_can_lehmann_fsm/_0397_ ;
 wire \heichips25_can_lehmann_fsm/_0398_ ;
 wire \heichips25_can_lehmann_fsm/_0399_ ;
 wire \heichips25_can_lehmann_fsm/_0400_ ;
 wire \heichips25_can_lehmann_fsm/_0401_ ;
 wire \heichips25_can_lehmann_fsm/_0402_ ;
 wire \heichips25_can_lehmann_fsm/_0403_ ;
 wire \heichips25_can_lehmann_fsm/_0404_ ;
 wire \heichips25_can_lehmann_fsm/_0405_ ;
 wire \heichips25_can_lehmann_fsm/_0406_ ;
 wire \heichips25_can_lehmann_fsm/_0407_ ;
 wire \heichips25_can_lehmann_fsm/_0408_ ;
 wire \heichips25_can_lehmann_fsm/_0409_ ;
 wire \heichips25_can_lehmann_fsm/_0410_ ;
 wire \heichips25_can_lehmann_fsm/_0411_ ;
 wire \heichips25_can_lehmann_fsm/_0412_ ;
 wire \heichips25_can_lehmann_fsm/_0413_ ;
 wire \heichips25_can_lehmann_fsm/_0414_ ;
 wire \heichips25_can_lehmann_fsm/_0415_ ;
 wire \heichips25_can_lehmann_fsm/_0416_ ;
 wire \heichips25_can_lehmann_fsm/_0417_ ;
 wire \heichips25_can_lehmann_fsm/_0418_ ;
 wire \heichips25_can_lehmann_fsm/_0419_ ;
 wire \heichips25_can_lehmann_fsm/_0420_ ;
 wire \heichips25_can_lehmann_fsm/_0421_ ;
 wire \heichips25_can_lehmann_fsm/_0422_ ;
 wire \heichips25_can_lehmann_fsm/_0423_ ;
 wire \heichips25_can_lehmann_fsm/_0424_ ;
 wire \heichips25_can_lehmann_fsm/_0425_ ;
 wire \heichips25_can_lehmann_fsm/_0426_ ;
 wire \heichips25_can_lehmann_fsm/_0427_ ;
 wire \heichips25_can_lehmann_fsm/_0428_ ;
 wire \heichips25_can_lehmann_fsm/_0429_ ;
 wire \heichips25_can_lehmann_fsm/_0430_ ;
 wire \heichips25_can_lehmann_fsm/_0431_ ;
 wire \heichips25_can_lehmann_fsm/_0432_ ;
 wire \heichips25_can_lehmann_fsm/_0433_ ;
 wire \heichips25_can_lehmann_fsm/_0434_ ;
 wire \heichips25_can_lehmann_fsm/_0435_ ;
 wire \heichips25_can_lehmann_fsm/_0436_ ;
 wire \heichips25_can_lehmann_fsm/_0437_ ;
 wire \heichips25_can_lehmann_fsm/_0438_ ;
 wire \heichips25_can_lehmann_fsm/_0439_ ;
 wire \heichips25_can_lehmann_fsm/_0440_ ;
 wire \heichips25_can_lehmann_fsm/_0441_ ;
 wire \heichips25_can_lehmann_fsm/_0442_ ;
 wire \heichips25_can_lehmann_fsm/_0443_ ;
 wire \heichips25_can_lehmann_fsm/_0444_ ;
 wire \heichips25_can_lehmann_fsm/_0445_ ;
 wire \heichips25_can_lehmann_fsm/_0446_ ;
 wire \heichips25_can_lehmann_fsm/_0447_ ;
 wire \heichips25_can_lehmann_fsm/_0448_ ;
 wire \heichips25_can_lehmann_fsm/_0449_ ;
 wire \heichips25_can_lehmann_fsm/_0450_ ;
 wire \heichips25_can_lehmann_fsm/_0451_ ;
 wire \heichips25_can_lehmann_fsm/_0452_ ;
 wire \heichips25_can_lehmann_fsm/_0453_ ;
 wire \heichips25_can_lehmann_fsm/_0454_ ;
 wire \heichips25_can_lehmann_fsm/_0455_ ;
 wire \heichips25_can_lehmann_fsm/_0456_ ;
 wire \heichips25_can_lehmann_fsm/_0457_ ;
 wire \heichips25_can_lehmann_fsm/_0458_ ;
 wire \heichips25_can_lehmann_fsm/_0459_ ;
 wire \heichips25_can_lehmann_fsm/_0460_ ;
 wire \heichips25_can_lehmann_fsm/_0461_ ;
 wire \heichips25_can_lehmann_fsm/_0462_ ;
 wire \heichips25_can_lehmann_fsm/_0463_ ;
 wire \heichips25_can_lehmann_fsm/_0464_ ;
 wire \heichips25_can_lehmann_fsm/_0465_ ;
 wire \heichips25_can_lehmann_fsm/_0466_ ;
 wire \heichips25_can_lehmann_fsm/_0467_ ;
 wire \heichips25_can_lehmann_fsm/_0468_ ;
 wire \heichips25_can_lehmann_fsm/_0469_ ;
 wire \heichips25_can_lehmann_fsm/_0470_ ;
 wire \heichips25_can_lehmann_fsm/_0471_ ;
 wire \heichips25_can_lehmann_fsm/_0472_ ;
 wire \heichips25_can_lehmann_fsm/_0473_ ;
 wire \heichips25_can_lehmann_fsm/_0474_ ;
 wire \heichips25_can_lehmann_fsm/_0475_ ;
 wire \heichips25_can_lehmann_fsm/_0476_ ;
 wire \heichips25_can_lehmann_fsm/_0477_ ;
 wire \heichips25_can_lehmann_fsm/_0478_ ;
 wire \heichips25_can_lehmann_fsm/_0479_ ;
 wire \heichips25_can_lehmann_fsm/_0480_ ;
 wire \heichips25_can_lehmann_fsm/_0481_ ;
 wire \heichips25_can_lehmann_fsm/_0482_ ;
 wire \heichips25_can_lehmann_fsm/_0483_ ;
 wire \heichips25_can_lehmann_fsm/_0484_ ;
 wire \heichips25_can_lehmann_fsm/_0485_ ;
 wire \heichips25_can_lehmann_fsm/_0486_ ;
 wire \heichips25_can_lehmann_fsm/_0487_ ;
 wire \heichips25_can_lehmann_fsm/_0488_ ;
 wire \heichips25_can_lehmann_fsm/_0489_ ;
 wire \heichips25_can_lehmann_fsm/_0490_ ;
 wire \heichips25_can_lehmann_fsm/_0491_ ;
 wire \heichips25_can_lehmann_fsm/_0492_ ;
 wire \heichips25_can_lehmann_fsm/_0493_ ;
 wire \heichips25_can_lehmann_fsm/_0494_ ;
 wire \heichips25_can_lehmann_fsm/_0495_ ;
 wire \heichips25_can_lehmann_fsm/_0496_ ;
 wire \heichips25_can_lehmann_fsm/_0497_ ;
 wire \heichips25_can_lehmann_fsm/_0498_ ;
 wire \heichips25_can_lehmann_fsm/_0499_ ;
 wire \heichips25_can_lehmann_fsm/_0500_ ;
 wire \heichips25_can_lehmann_fsm/_0501_ ;
 wire \heichips25_can_lehmann_fsm/_0502_ ;
 wire \heichips25_can_lehmann_fsm/_0503_ ;
 wire \heichips25_can_lehmann_fsm/_0504_ ;
 wire \heichips25_can_lehmann_fsm/_0505_ ;
 wire \heichips25_can_lehmann_fsm/_0506_ ;
 wire \heichips25_can_lehmann_fsm/_0507_ ;
 wire \heichips25_can_lehmann_fsm/_0508_ ;
 wire \heichips25_can_lehmann_fsm/_0509_ ;
 wire \heichips25_can_lehmann_fsm/_0510_ ;
 wire \heichips25_can_lehmann_fsm/_0511_ ;
 wire \heichips25_can_lehmann_fsm/_0512_ ;
 wire \heichips25_can_lehmann_fsm/_0513_ ;
 wire \heichips25_can_lehmann_fsm/_0514_ ;
 wire \heichips25_can_lehmann_fsm/_0515_ ;
 wire \heichips25_can_lehmann_fsm/_0516_ ;
 wire \heichips25_can_lehmann_fsm/_0517_ ;
 wire \heichips25_can_lehmann_fsm/_0518_ ;
 wire \heichips25_can_lehmann_fsm/_0519_ ;
 wire \heichips25_can_lehmann_fsm/_0520_ ;
 wire \heichips25_can_lehmann_fsm/_0521_ ;
 wire \heichips25_can_lehmann_fsm/_0522_ ;
 wire \heichips25_can_lehmann_fsm/_0523_ ;
 wire \heichips25_can_lehmann_fsm/_0524_ ;
 wire \heichips25_can_lehmann_fsm/_0525_ ;
 wire \heichips25_can_lehmann_fsm/_0526_ ;
 wire \heichips25_can_lehmann_fsm/_0527_ ;
 wire \heichips25_can_lehmann_fsm/_0528_ ;
 wire \heichips25_can_lehmann_fsm/_0529_ ;
 wire \heichips25_can_lehmann_fsm/_0530_ ;
 wire \heichips25_can_lehmann_fsm/_0531_ ;
 wire \heichips25_can_lehmann_fsm/_0532_ ;
 wire \heichips25_can_lehmann_fsm/_0533_ ;
 wire \heichips25_can_lehmann_fsm/_0534_ ;
 wire \heichips25_can_lehmann_fsm/_0535_ ;
 wire \heichips25_can_lehmann_fsm/_0536_ ;
 wire \heichips25_can_lehmann_fsm/_0537_ ;
 wire \heichips25_can_lehmann_fsm/_0538_ ;
 wire \heichips25_can_lehmann_fsm/_0539_ ;
 wire \heichips25_can_lehmann_fsm/_0540_ ;
 wire \heichips25_can_lehmann_fsm/_0541_ ;
 wire \heichips25_can_lehmann_fsm/_0542_ ;
 wire \heichips25_can_lehmann_fsm/_0543_ ;
 wire \heichips25_can_lehmann_fsm/_0544_ ;
 wire \heichips25_can_lehmann_fsm/_0545_ ;
 wire \heichips25_can_lehmann_fsm/_0546_ ;
 wire \heichips25_can_lehmann_fsm/_0547_ ;
 wire \heichips25_can_lehmann_fsm/_0548_ ;
 wire \heichips25_can_lehmann_fsm/_0549_ ;
 wire \heichips25_can_lehmann_fsm/_0550_ ;
 wire \heichips25_can_lehmann_fsm/_0551_ ;
 wire \heichips25_can_lehmann_fsm/_0552_ ;
 wire \heichips25_can_lehmann_fsm/_0553_ ;
 wire \heichips25_can_lehmann_fsm/_0554_ ;
 wire \heichips25_can_lehmann_fsm/_0555_ ;
 wire \heichips25_can_lehmann_fsm/_0556_ ;
 wire \heichips25_can_lehmann_fsm/_0557_ ;
 wire \heichips25_can_lehmann_fsm/_0558_ ;
 wire \heichips25_can_lehmann_fsm/_0559_ ;
 wire \heichips25_can_lehmann_fsm/_0560_ ;
 wire \heichips25_can_lehmann_fsm/_0561_ ;
 wire \heichips25_can_lehmann_fsm/_0562_ ;
 wire \heichips25_can_lehmann_fsm/_0563_ ;
 wire \heichips25_can_lehmann_fsm/_0564_ ;
 wire \heichips25_can_lehmann_fsm/_0565_ ;
 wire \heichips25_can_lehmann_fsm/_0566_ ;
 wire \heichips25_can_lehmann_fsm/_0567_ ;
 wire \heichips25_can_lehmann_fsm/_0568_ ;
 wire \heichips25_can_lehmann_fsm/_0569_ ;
 wire \heichips25_can_lehmann_fsm/_0570_ ;
 wire \heichips25_can_lehmann_fsm/_0571_ ;
 wire \heichips25_can_lehmann_fsm/_0572_ ;
 wire \heichips25_can_lehmann_fsm/_0573_ ;
 wire \heichips25_can_lehmann_fsm/_0574_ ;
 wire \heichips25_can_lehmann_fsm/_0575_ ;
 wire \heichips25_can_lehmann_fsm/_0576_ ;
 wire \heichips25_can_lehmann_fsm/_0577_ ;
 wire \heichips25_can_lehmann_fsm/_0578_ ;
 wire \heichips25_can_lehmann_fsm/_0579_ ;
 wire \heichips25_can_lehmann_fsm/_0580_ ;
 wire \heichips25_can_lehmann_fsm/_0581_ ;
 wire \heichips25_can_lehmann_fsm/_0582_ ;
 wire \heichips25_can_lehmann_fsm/_0583_ ;
 wire \heichips25_can_lehmann_fsm/_0584_ ;
 wire \heichips25_can_lehmann_fsm/_0585_ ;
 wire \heichips25_can_lehmann_fsm/_0586_ ;
 wire \heichips25_can_lehmann_fsm/_0587_ ;
 wire \heichips25_can_lehmann_fsm/_0588_ ;
 wire \heichips25_can_lehmann_fsm/_0589_ ;
 wire \heichips25_can_lehmann_fsm/_0590_ ;
 wire \heichips25_can_lehmann_fsm/_0591_ ;
 wire \heichips25_can_lehmann_fsm/_0592_ ;
 wire \heichips25_can_lehmann_fsm/_0593_ ;
 wire \heichips25_can_lehmann_fsm/_0594_ ;
 wire \heichips25_can_lehmann_fsm/_0595_ ;
 wire \heichips25_can_lehmann_fsm/_0596_ ;
 wire \heichips25_can_lehmann_fsm/_0597_ ;
 wire \heichips25_can_lehmann_fsm/_0598_ ;
 wire \heichips25_can_lehmann_fsm/_0599_ ;
 wire \heichips25_can_lehmann_fsm/_0600_ ;
 wire \heichips25_can_lehmann_fsm/_0601_ ;
 wire \heichips25_can_lehmann_fsm/_0602_ ;
 wire \heichips25_can_lehmann_fsm/_0603_ ;
 wire \heichips25_can_lehmann_fsm/_0604_ ;
 wire \heichips25_can_lehmann_fsm/_0605_ ;
 wire \heichips25_can_lehmann_fsm/_0606_ ;
 wire \heichips25_can_lehmann_fsm/_0607_ ;
 wire \heichips25_can_lehmann_fsm/_0608_ ;
 wire \heichips25_can_lehmann_fsm/_0609_ ;
 wire \heichips25_can_lehmann_fsm/_0610_ ;
 wire \heichips25_can_lehmann_fsm/_0611_ ;
 wire \heichips25_can_lehmann_fsm/_0612_ ;
 wire \heichips25_can_lehmann_fsm/_0613_ ;
 wire \heichips25_can_lehmann_fsm/_0614_ ;
 wire \heichips25_can_lehmann_fsm/_0615_ ;
 wire \heichips25_can_lehmann_fsm/_0616_ ;
 wire \heichips25_can_lehmann_fsm/_0617_ ;
 wire \heichips25_can_lehmann_fsm/_0618_ ;
 wire \heichips25_can_lehmann_fsm/_0619_ ;
 wire \heichips25_can_lehmann_fsm/_0620_ ;
 wire \heichips25_can_lehmann_fsm/_0621_ ;
 wire \heichips25_can_lehmann_fsm/_0622_ ;
 wire \heichips25_can_lehmann_fsm/_0623_ ;
 wire \heichips25_can_lehmann_fsm/_0624_ ;
 wire \heichips25_can_lehmann_fsm/_0625_ ;
 wire \heichips25_can_lehmann_fsm/_0626_ ;
 wire \heichips25_can_lehmann_fsm/_0627_ ;
 wire \heichips25_can_lehmann_fsm/_0628_ ;
 wire \heichips25_can_lehmann_fsm/_0629_ ;
 wire \heichips25_can_lehmann_fsm/_0630_ ;
 wire \heichips25_can_lehmann_fsm/_0631_ ;
 wire \heichips25_can_lehmann_fsm/_0632_ ;
 wire \heichips25_can_lehmann_fsm/_0633_ ;
 wire \heichips25_can_lehmann_fsm/_0634_ ;
 wire \heichips25_can_lehmann_fsm/_0635_ ;
 wire \heichips25_can_lehmann_fsm/_0636_ ;
 wire \heichips25_can_lehmann_fsm/_0637_ ;
 wire \heichips25_can_lehmann_fsm/_0638_ ;
 wire \heichips25_can_lehmann_fsm/_0639_ ;
 wire \heichips25_can_lehmann_fsm/_0640_ ;
 wire \heichips25_can_lehmann_fsm/_0641_ ;
 wire \heichips25_can_lehmann_fsm/_0642_ ;
 wire \heichips25_can_lehmann_fsm/_0643_ ;
 wire \heichips25_can_lehmann_fsm/_0644_ ;
 wire \heichips25_can_lehmann_fsm/_0645_ ;
 wire \heichips25_can_lehmann_fsm/_0646_ ;
 wire \heichips25_can_lehmann_fsm/_0647_ ;
 wire \heichips25_can_lehmann_fsm/_0648_ ;
 wire \heichips25_can_lehmann_fsm/_0649_ ;
 wire \heichips25_can_lehmann_fsm/_0650_ ;
 wire \heichips25_can_lehmann_fsm/_0651_ ;
 wire \heichips25_can_lehmann_fsm/_0652_ ;
 wire \heichips25_can_lehmann_fsm/_0653_ ;
 wire \heichips25_can_lehmann_fsm/_0654_ ;
 wire \heichips25_can_lehmann_fsm/_0655_ ;
 wire \heichips25_can_lehmann_fsm/_0656_ ;
 wire \heichips25_can_lehmann_fsm/_0657_ ;
 wire \heichips25_can_lehmann_fsm/_0658_ ;
 wire \heichips25_can_lehmann_fsm/_0659_ ;
 wire \heichips25_can_lehmann_fsm/_0660_ ;
 wire \heichips25_can_lehmann_fsm/_0661_ ;
 wire \heichips25_can_lehmann_fsm/_0662_ ;
 wire \heichips25_can_lehmann_fsm/_0663_ ;
 wire \heichips25_can_lehmann_fsm/_0664_ ;
 wire \heichips25_can_lehmann_fsm/_0665_ ;
 wire \heichips25_can_lehmann_fsm/_0666_ ;
 wire \heichips25_can_lehmann_fsm/_0667_ ;
 wire \heichips25_can_lehmann_fsm/_0668_ ;
 wire \heichips25_can_lehmann_fsm/_0669_ ;
 wire \heichips25_can_lehmann_fsm/_0670_ ;
 wire \heichips25_can_lehmann_fsm/_0671_ ;
 wire \heichips25_can_lehmann_fsm/_0672_ ;
 wire \heichips25_can_lehmann_fsm/_0673_ ;
 wire \heichips25_can_lehmann_fsm/_0674_ ;
 wire \heichips25_can_lehmann_fsm/_0675_ ;
 wire \heichips25_can_lehmann_fsm/_0676_ ;
 wire \heichips25_can_lehmann_fsm/_0677_ ;
 wire \heichips25_can_lehmann_fsm/_0678_ ;
 wire \heichips25_can_lehmann_fsm/_0679_ ;
 wire \heichips25_can_lehmann_fsm/_0680_ ;
 wire \heichips25_can_lehmann_fsm/_0681_ ;
 wire \heichips25_can_lehmann_fsm/_0682_ ;
 wire \heichips25_can_lehmann_fsm/_0683_ ;
 wire \heichips25_can_lehmann_fsm/_0684_ ;
 wire \heichips25_can_lehmann_fsm/_0685_ ;
 wire \heichips25_can_lehmann_fsm/_0686_ ;
 wire \heichips25_can_lehmann_fsm/_0687_ ;
 wire \heichips25_can_lehmann_fsm/_0688_ ;
 wire \heichips25_can_lehmann_fsm/_0689_ ;
 wire \heichips25_can_lehmann_fsm/_0690_ ;
 wire \heichips25_can_lehmann_fsm/_0691_ ;
 wire \heichips25_can_lehmann_fsm/_0692_ ;
 wire \heichips25_can_lehmann_fsm/_0693_ ;
 wire \heichips25_can_lehmann_fsm/_0694_ ;
 wire \heichips25_can_lehmann_fsm/_0695_ ;
 wire \heichips25_can_lehmann_fsm/_0696_ ;
 wire \heichips25_can_lehmann_fsm/_0697_ ;
 wire \heichips25_can_lehmann_fsm/_0698_ ;
 wire \heichips25_can_lehmann_fsm/_0699_ ;
 wire \heichips25_can_lehmann_fsm/_0700_ ;
 wire \heichips25_can_lehmann_fsm/_0701_ ;
 wire \heichips25_can_lehmann_fsm/_0702_ ;
 wire \heichips25_can_lehmann_fsm/_0703_ ;
 wire \heichips25_can_lehmann_fsm/_0704_ ;
 wire \heichips25_can_lehmann_fsm/_0705_ ;
 wire \heichips25_can_lehmann_fsm/_0706_ ;
 wire \heichips25_can_lehmann_fsm/_0707_ ;
 wire \heichips25_can_lehmann_fsm/_0708_ ;
 wire \heichips25_can_lehmann_fsm/_0709_ ;
 wire \heichips25_can_lehmann_fsm/_0710_ ;
 wire \heichips25_can_lehmann_fsm/_0711_ ;
 wire \heichips25_can_lehmann_fsm/_0712_ ;
 wire \heichips25_can_lehmann_fsm/_0713_ ;
 wire \heichips25_can_lehmann_fsm/_0714_ ;
 wire \heichips25_can_lehmann_fsm/_0715_ ;
 wire \heichips25_can_lehmann_fsm/_0716_ ;
 wire \heichips25_can_lehmann_fsm/_0717_ ;
 wire \heichips25_can_lehmann_fsm/_0718_ ;
 wire \heichips25_can_lehmann_fsm/_0719_ ;
 wire \heichips25_can_lehmann_fsm/_0720_ ;
 wire \heichips25_can_lehmann_fsm/_0721_ ;
 wire \heichips25_can_lehmann_fsm/_0722_ ;
 wire \heichips25_can_lehmann_fsm/_0723_ ;
 wire \heichips25_can_lehmann_fsm/_0724_ ;
 wire \heichips25_can_lehmann_fsm/_0725_ ;
 wire \heichips25_can_lehmann_fsm/_0726_ ;
 wire \heichips25_can_lehmann_fsm/_0727_ ;
 wire \heichips25_can_lehmann_fsm/_0728_ ;
 wire \heichips25_can_lehmann_fsm/_0729_ ;
 wire \heichips25_can_lehmann_fsm/_0730_ ;
 wire \heichips25_can_lehmann_fsm/_0731_ ;
 wire \heichips25_can_lehmann_fsm/_0732_ ;
 wire \heichips25_can_lehmann_fsm/_0733_ ;
 wire \heichips25_can_lehmann_fsm/_0734_ ;
 wire \heichips25_can_lehmann_fsm/_0735_ ;
 wire \heichips25_can_lehmann_fsm/_0736_ ;
 wire \heichips25_can_lehmann_fsm/_0737_ ;
 wire \heichips25_can_lehmann_fsm/_0738_ ;
 wire \heichips25_can_lehmann_fsm/_0739_ ;
 wire \heichips25_can_lehmann_fsm/_0740_ ;
 wire \heichips25_can_lehmann_fsm/_0741_ ;
 wire \heichips25_can_lehmann_fsm/_0742_ ;
 wire \heichips25_can_lehmann_fsm/_0743_ ;
 wire \heichips25_can_lehmann_fsm/_0744_ ;
 wire \heichips25_can_lehmann_fsm/_0745_ ;
 wire \heichips25_can_lehmann_fsm/_0746_ ;
 wire \heichips25_can_lehmann_fsm/_0747_ ;
 wire \heichips25_can_lehmann_fsm/_0748_ ;
 wire \heichips25_can_lehmann_fsm/_0749_ ;
 wire \heichips25_can_lehmann_fsm/_0750_ ;
 wire \heichips25_can_lehmann_fsm/_0751_ ;
 wire \heichips25_can_lehmann_fsm/_0752_ ;
 wire \heichips25_can_lehmann_fsm/_0753_ ;
 wire \heichips25_can_lehmann_fsm/_0754_ ;
 wire \heichips25_can_lehmann_fsm/_0755_ ;
 wire \heichips25_can_lehmann_fsm/_0756_ ;
 wire \heichips25_can_lehmann_fsm/_0757_ ;
 wire \heichips25_can_lehmann_fsm/_0758_ ;
 wire \heichips25_can_lehmann_fsm/_0759_ ;
 wire \heichips25_can_lehmann_fsm/_0760_ ;
 wire \heichips25_can_lehmann_fsm/_0761_ ;
 wire \heichips25_can_lehmann_fsm/_0762_ ;
 wire \heichips25_can_lehmann_fsm/_0763_ ;
 wire \heichips25_can_lehmann_fsm/_0764_ ;
 wire \heichips25_can_lehmann_fsm/_0765_ ;
 wire \heichips25_can_lehmann_fsm/_0766_ ;
 wire \heichips25_can_lehmann_fsm/_0767_ ;
 wire \heichips25_can_lehmann_fsm/_0768_ ;
 wire \heichips25_can_lehmann_fsm/_0769_ ;
 wire \heichips25_can_lehmann_fsm/_0770_ ;
 wire \heichips25_can_lehmann_fsm/_0771_ ;
 wire \heichips25_can_lehmann_fsm/_0772_ ;
 wire \heichips25_can_lehmann_fsm/_0773_ ;
 wire \heichips25_can_lehmann_fsm/_0774_ ;
 wire \heichips25_can_lehmann_fsm/_0775_ ;
 wire \heichips25_can_lehmann_fsm/_0776_ ;
 wire \heichips25_can_lehmann_fsm/_0777_ ;
 wire \heichips25_can_lehmann_fsm/_0778_ ;
 wire \heichips25_can_lehmann_fsm/_0779_ ;
 wire \heichips25_can_lehmann_fsm/_0780_ ;
 wire \heichips25_can_lehmann_fsm/_0781_ ;
 wire \heichips25_can_lehmann_fsm/_0782_ ;
 wire \heichips25_can_lehmann_fsm/_0783_ ;
 wire \heichips25_can_lehmann_fsm/_0784_ ;
 wire \heichips25_can_lehmann_fsm/_0785_ ;
 wire \heichips25_can_lehmann_fsm/_0786_ ;
 wire \heichips25_can_lehmann_fsm/_0787_ ;
 wire \heichips25_can_lehmann_fsm/_0788_ ;
 wire \heichips25_can_lehmann_fsm/_0789_ ;
 wire \heichips25_can_lehmann_fsm/_0790_ ;
 wire \heichips25_can_lehmann_fsm/_0791_ ;
 wire \heichips25_can_lehmann_fsm/_0792_ ;
 wire \heichips25_can_lehmann_fsm/_0793_ ;
 wire \heichips25_can_lehmann_fsm/_0794_ ;
 wire \heichips25_can_lehmann_fsm/_0795_ ;
 wire \heichips25_can_lehmann_fsm/_0796_ ;
 wire \heichips25_can_lehmann_fsm/_0797_ ;
 wire \heichips25_can_lehmann_fsm/_0798_ ;
 wire \heichips25_can_lehmann_fsm/_0799_ ;
 wire \heichips25_can_lehmann_fsm/_0800_ ;
 wire \heichips25_can_lehmann_fsm/_0801_ ;
 wire \heichips25_can_lehmann_fsm/_0802_ ;
 wire \heichips25_can_lehmann_fsm/_0803_ ;
 wire \heichips25_can_lehmann_fsm/_0804_ ;
 wire \heichips25_can_lehmann_fsm/_0805_ ;
 wire \heichips25_can_lehmann_fsm/_0806_ ;
 wire \heichips25_can_lehmann_fsm/_0807_ ;
 wire \heichips25_can_lehmann_fsm/_0808_ ;
 wire \heichips25_can_lehmann_fsm/_0809_ ;
 wire \heichips25_can_lehmann_fsm/_0810_ ;
 wire \heichips25_can_lehmann_fsm/_0811_ ;
 wire \heichips25_can_lehmann_fsm/_0812_ ;
 wire \heichips25_can_lehmann_fsm/_0813_ ;
 wire \heichips25_can_lehmann_fsm/_0814_ ;
 wire \heichips25_can_lehmann_fsm/_0815_ ;
 wire \heichips25_can_lehmann_fsm/_0816_ ;
 wire \heichips25_can_lehmann_fsm/_0817_ ;
 wire \heichips25_can_lehmann_fsm/_0818_ ;
 wire \heichips25_can_lehmann_fsm/_0819_ ;
 wire \heichips25_can_lehmann_fsm/_0820_ ;
 wire \heichips25_can_lehmann_fsm/_0821_ ;
 wire \heichips25_can_lehmann_fsm/_0822_ ;
 wire \heichips25_can_lehmann_fsm/_0823_ ;
 wire \heichips25_can_lehmann_fsm/_0824_ ;
 wire \heichips25_can_lehmann_fsm/_0825_ ;
 wire \heichips25_can_lehmann_fsm/_0826_ ;
 wire \heichips25_can_lehmann_fsm/_0827_ ;
 wire \heichips25_can_lehmann_fsm/_0828_ ;
 wire \heichips25_can_lehmann_fsm/_0829_ ;
 wire \heichips25_can_lehmann_fsm/_0830_ ;
 wire \heichips25_can_lehmann_fsm/_0831_ ;
 wire \heichips25_can_lehmann_fsm/_0832_ ;
 wire \heichips25_can_lehmann_fsm/_0833_ ;
 wire \heichips25_can_lehmann_fsm/_0834_ ;
 wire \heichips25_can_lehmann_fsm/_0835_ ;
 wire \heichips25_can_lehmann_fsm/_0836_ ;
 wire \heichips25_can_lehmann_fsm/_0837_ ;
 wire \heichips25_can_lehmann_fsm/_0838_ ;
 wire \heichips25_can_lehmann_fsm/_0839_ ;
 wire \heichips25_can_lehmann_fsm/_0840_ ;
 wire \heichips25_can_lehmann_fsm/_0841_ ;
 wire \heichips25_can_lehmann_fsm/_0842_ ;
 wire \heichips25_can_lehmann_fsm/_0843_ ;
 wire \heichips25_can_lehmann_fsm/_0844_ ;
 wire \heichips25_can_lehmann_fsm/_0845_ ;
 wire \heichips25_can_lehmann_fsm/_0846_ ;
 wire \heichips25_can_lehmann_fsm/_0847_ ;
 wire \heichips25_can_lehmann_fsm/_0848_ ;
 wire \heichips25_can_lehmann_fsm/_0849_ ;
 wire \heichips25_can_lehmann_fsm/_0850_ ;
 wire \heichips25_can_lehmann_fsm/_0851_ ;
 wire \heichips25_can_lehmann_fsm/_0852_ ;
 wire \heichips25_can_lehmann_fsm/_0853_ ;
 wire \heichips25_can_lehmann_fsm/_0854_ ;
 wire \heichips25_can_lehmann_fsm/_0855_ ;
 wire \heichips25_can_lehmann_fsm/_0856_ ;
 wire \heichips25_can_lehmann_fsm/_0857_ ;
 wire \heichips25_can_lehmann_fsm/_0858_ ;
 wire \heichips25_can_lehmann_fsm/_0859_ ;
 wire \heichips25_can_lehmann_fsm/_0860_ ;
 wire \heichips25_can_lehmann_fsm/_0861_ ;
 wire \heichips25_can_lehmann_fsm/_0862_ ;
 wire \heichips25_can_lehmann_fsm/_0863_ ;
 wire \heichips25_can_lehmann_fsm/_0864_ ;
 wire \heichips25_can_lehmann_fsm/_0865_ ;
 wire \heichips25_can_lehmann_fsm/_0866_ ;
 wire \heichips25_can_lehmann_fsm/_0867_ ;
 wire \heichips25_can_lehmann_fsm/_0868_ ;
 wire \heichips25_can_lehmann_fsm/_0869_ ;
 wire \heichips25_can_lehmann_fsm/_0870_ ;
 wire \heichips25_can_lehmann_fsm/_0871_ ;
 wire \heichips25_can_lehmann_fsm/_0872_ ;
 wire \heichips25_can_lehmann_fsm/_0873_ ;
 wire \heichips25_can_lehmann_fsm/_0874_ ;
 wire \heichips25_can_lehmann_fsm/_0875_ ;
 wire \heichips25_can_lehmann_fsm/_0876_ ;
 wire \heichips25_can_lehmann_fsm/_0877_ ;
 wire \heichips25_can_lehmann_fsm/_0878_ ;
 wire \heichips25_can_lehmann_fsm/_0879_ ;
 wire \heichips25_can_lehmann_fsm/_0880_ ;
 wire \heichips25_can_lehmann_fsm/_0881_ ;
 wire \heichips25_can_lehmann_fsm/_0882_ ;
 wire \heichips25_can_lehmann_fsm/_0883_ ;
 wire \heichips25_can_lehmann_fsm/_0884_ ;
 wire \heichips25_can_lehmann_fsm/_0885_ ;
 wire \heichips25_can_lehmann_fsm/_0886_ ;
 wire \heichips25_can_lehmann_fsm/_0887_ ;
 wire \heichips25_can_lehmann_fsm/_0888_ ;
 wire \heichips25_can_lehmann_fsm/_0889_ ;
 wire \heichips25_can_lehmann_fsm/_0890_ ;
 wire \heichips25_can_lehmann_fsm/_0891_ ;
 wire \heichips25_can_lehmann_fsm/_0892_ ;
 wire \heichips25_can_lehmann_fsm/_0893_ ;
 wire \heichips25_can_lehmann_fsm/_0894_ ;
 wire \heichips25_can_lehmann_fsm/_0895_ ;
 wire \heichips25_can_lehmann_fsm/_0896_ ;
 wire \heichips25_can_lehmann_fsm/_0897_ ;
 wire \heichips25_can_lehmann_fsm/_0898_ ;
 wire \heichips25_can_lehmann_fsm/_0899_ ;
 wire \heichips25_can_lehmann_fsm/_0900_ ;
 wire \heichips25_can_lehmann_fsm/_0901_ ;
 wire \heichips25_can_lehmann_fsm/_0902_ ;
 wire \heichips25_can_lehmann_fsm/_0903_ ;
 wire \heichips25_can_lehmann_fsm/_0904_ ;
 wire \heichips25_can_lehmann_fsm/_0905_ ;
 wire \heichips25_can_lehmann_fsm/_0906_ ;
 wire \heichips25_can_lehmann_fsm/_0907_ ;
 wire \heichips25_can_lehmann_fsm/_0908_ ;
 wire \heichips25_can_lehmann_fsm/_0909_ ;
 wire \heichips25_can_lehmann_fsm/_0910_ ;
 wire \heichips25_can_lehmann_fsm/_0911_ ;
 wire \heichips25_can_lehmann_fsm/_0912_ ;
 wire \heichips25_can_lehmann_fsm/_0913_ ;
 wire \heichips25_can_lehmann_fsm/_0914_ ;
 wire \heichips25_can_lehmann_fsm/_0915_ ;
 wire \heichips25_can_lehmann_fsm/_0916_ ;
 wire \heichips25_can_lehmann_fsm/_0917_ ;
 wire \heichips25_can_lehmann_fsm/_0918_ ;
 wire \heichips25_can_lehmann_fsm/_0919_ ;
 wire \heichips25_can_lehmann_fsm/_0920_ ;
 wire \heichips25_can_lehmann_fsm/_0921_ ;
 wire \heichips25_can_lehmann_fsm/_0922_ ;
 wire \heichips25_can_lehmann_fsm/_0923_ ;
 wire \heichips25_can_lehmann_fsm/_0924_ ;
 wire \heichips25_can_lehmann_fsm/_0925_ ;
 wire \heichips25_can_lehmann_fsm/_0926_ ;
 wire \heichips25_can_lehmann_fsm/_0927_ ;
 wire \heichips25_can_lehmann_fsm/_0928_ ;
 wire \heichips25_can_lehmann_fsm/_0929_ ;
 wire \heichips25_can_lehmann_fsm/_0930_ ;
 wire \heichips25_can_lehmann_fsm/_0931_ ;
 wire \heichips25_can_lehmann_fsm/_0932_ ;
 wire \heichips25_can_lehmann_fsm/_0933_ ;
 wire \heichips25_can_lehmann_fsm/_0934_ ;
 wire \heichips25_can_lehmann_fsm/_0935_ ;
 wire \heichips25_can_lehmann_fsm/_0936_ ;
 wire \heichips25_can_lehmann_fsm/_0937_ ;
 wire \heichips25_can_lehmann_fsm/_0938_ ;
 wire \heichips25_can_lehmann_fsm/_0939_ ;
 wire \heichips25_can_lehmann_fsm/_0940_ ;
 wire \heichips25_can_lehmann_fsm/_0941_ ;
 wire \heichips25_can_lehmann_fsm/_0942_ ;
 wire \heichips25_can_lehmann_fsm/_0943_ ;
 wire \heichips25_can_lehmann_fsm/_0944_ ;
 wire \heichips25_can_lehmann_fsm/_0945_ ;
 wire \heichips25_can_lehmann_fsm/_0946_ ;
 wire \heichips25_can_lehmann_fsm/_0947_ ;
 wire \heichips25_can_lehmann_fsm/_0948_ ;
 wire \heichips25_can_lehmann_fsm/_0949_ ;
 wire \heichips25_can_lehmann_fsm/_0950_ ;
 wire \heichips25_can_lehmann_fsm/_0951_ ;
 wire \heichips25_can_lehmann_fsm/_0952_ ;
 wire \heichips25_can_lehmann_fsm/_0953_ ;
 wire \heichips25_can_lehmann_fsm/_0954_ ;
 wire \heichips25_can_lehmann_fsm/_0955_ ;
 wire \heichips25_can_lehmann_fsm/_0956_ ;
 wire \heichips25_can_lehmann_fsm/_0957_ ;
 wire \heichips25_can_lehmann_fsm/_0958_ ;
 wire \heichips25_can_lehmann_fsm/_0959_ ;
 wire \heichips25_can_lehmann_fsm/_0960_ ;
 wire \heichips25_can_lehmann_fsm/_0961_ ;
 wire \heichips25_can_lehmann_fsm/_0962_ ;
 wire \heichips25_can_lehmann_fsm/_0963_ ;
 wire \heichips25_can_lehmann_fsm/_0964_ ;
 wire \heichips25_can_lehmann_fsm/_0965_ ;
 wire \heichips25_can_lehmann_fsm/_0966_ ;
 wire \heichips25_can_lehmann_fsm/_0967_ ;
 wire \heichips25_can_lehmann_fsm/_0968_ ;
 wire \heichips25_can_lehmann_fsm/_0969_ ;
 wire \heichips25_can_lehmann_fsm/_0970_ ;
 wire \heichips25_can_lehmann_fsm/_0971_ ;
 wire \heichips25_can_lehmann_fsm/_0972_ ;
 wire \heichips25_can_lehmann_fsm/_0973_ ;
 wire \heichips25_can_lehmann_fsm/_0974_ ;
 wire \heichips25_can_lehmann_fsm/_0975_ ;
 wire \heichips25_can_lehmann_fsm/_0976_ ;
 wire \heichips25_can_lehmann_fsm/_0977_ ;
 wire \heichips25_can_lehmann_fsm/_0978_ ;
 wire \heichips25_can_lehmann_fsm/_0979_ ;
 wire \heichips25_can_lehmann_fsm/_0980_ ;
 wire \heichips25_can_lehmann_fsm/_0981_ ;
 wire \heichips25_can_lehmann_fsm/_0982_ ;
 wire \heichips25_can_lehmann_fsm/_0983_ ;
 wire \heichips25_can_lehmann_fsm/_0984_ ;
 wire \heichips25_can_lehmann_fsm/_0985_ ;
 wire \heichips25_can_lehmann_fsm/_0986_ ;
 wire \heichips25_can_lehmann_fsm/_0987_ ;
 wire \heichips25_can_lehmann_fsm/_0988_ ;
 wire \heichips25_can_lehmann_fsm/_0989_ ;
 wire \heichips25_can_lehmann_fsm/_0990_ ;
 wire \heichips25_can_lehmann_fsm/_0991_ ;
 wire \heichips25_can_lehmann_fsm/_0992_ ;
 wire \heichips25_can_lehmann_fsm/_0993_ ;
 wire \heichips25_can_lehmann_fsm/_0994_ ;
 wire \heichips25_can_lehmann_fsm/_0995_ ;
 wire \heichips25_can_lehmann_fsm/_0996_ ;
 wire \heichips25_can_lehmann_fsm/_0997_ ;
 wire \heichips25_can_lehmann_fsm/_0998_ ;
 wire \heichips25_can_lehmann_fsm/_0999_ ;
 wire \heichips25_can_lehmann_fsm/_1000_ ;
 wire \heichips25_can_lehmann_fsm/_1001_ ;
 wire \heichips25_can_lehmann_fsm/_1002_ ;
 wire \heichips25_can_lehmann_fsm/_1003_ ;
 wire \heichips25_can_lehmann_fsm/_1004_ ;
 wire \heichips25_can_lehmann_fsm/_1005_ ;
 wire \heichips25_can_lehmann_fsm/_1006_ ;
 wire \heichips25_can_lehmann_fsm/_1007_ ;
 wire \heichips25_can_lehmann_fsm/_1008_ ;
 wire \heichips25_can_lehmann_fsm/_1009_ ;
 wire \heichips25_can_lehmann_fsm/_1010_ ;
 wire \heichips25_can_lehmann_fsm/_1011_ ;
 wire \heichips25_can_lehmann_fsm/_1012_ ;
 wire \heichips25_can_lehmann_fsm/_1013_ ;
 wire \heichips25_can_lehmann_fsm/_1014_ ;
 wire \heichips25_can_lehmann_fsm/_1015_ ;
 wire \heichips25_can_lehmann_fsm/_1016_ ;
 wire \heichips25_can_lehmann_fsm/_1017_ ;
 wire \heichips25_can_lehmann_fsm/_1018_ ;
 wire \heichips25_can_lehmann_fsm/_1019_ ;
 wire \heichips25_can_lehmann_fsm/_1020_ ;
 wire \heichips25_can_lehmann_fsm/_1021_ ;
 wire \heichips25_can_lehmann_fsm/_1022_ ;
 wire \heichips25_can_lehmann_fsm/_1023_ ;
 wire \heichips25_can_lehmann_fsm/_1024_ ;
 wire \heichips25_can_lehmann_fsm/_1025_ ;
 wire \heichips25_can_lehmann_fsm/_1026_ ;
 wire \heichips25_can_lehmann_fsm/_1027_ ;
 wire \heichips25_can_lehmann_fsm/_1028_ ;
 wire \heichips25_can_lehmann_fsm/_1029_ ;
 wire \heichips25_can_lehmann_fsm/_1030_ ;
 wire \heichips25_can_lehmann_fsm/_1031_ ;
 wire \heichips25_can_lehmann_fsm/_1032_ ;
 wire \heichips25_can_lehmann_fsm/_1033_ ;
 wire \heichips25_can_lehmann_fsm/_1034_ ;
 wire \heichips25_can_lehmann_fsm/_1035_ ;
 wire \heichips25_can_lehmann_fsm/_1036_ ;
 wire \heichips25_can_lehmann_fsm/_1037_ ;
 wire \heichips25_can_lehmann_fsm/_1038_ ;
 wire \heichips25_can_lehmann_fsm/_1039_ ;
 wire \heichips25_can_lehmann_fsm/_1040_ ;
 wire \heichips25_can_lehmann_fsm/_1041_ ;
 wire \heichips25_can_lehmann_fsm/_1042_ ;
 wire \heichips25_can_lehmann_fsm/_1043_ ;
 wire \heichips25_can_lehmann_fsm/_1044_ ;
 wire \heichips25_can_lehmann_fsm/_1045_ ;
 wire \heichips25_can_lehmann_fsm/_1046_ ;
 wire \heichips25_can_lehmann_fsm/_1047_ ;
 wire \heichips25_can_lehmann_fsm/_1048_ ;
 wire \heichips25_can_lehmann_fsm/_1049_ ;
 wire \heichips25_can_lehmann_fsm/_1050_ ;
 wire \heichips25_can_lehmann_fsm/_1051_ ;
 wire \heichips25_can_lehmann_fsm/_1052_ ;
 wire \heichips25_can_lehmann_fsm/_1053_ ;
 wire \heichips25_can_lehmann_fsm/_1054_ ;
 wire \heichips25_can_lehmann_fsm/_1055_ ;
 wire \heichips25_can_lehmann_fsm/_1056_ ;
 wire \heichips25_can_lehmann_fsm/_1057_ ;
 wire \heichips25_can_lehmann_fsm/_1058_ ;
 wire \heichips25_can_lehmann_fsm/_1059_ ;
 wire \heichips25_can_lehmann_fsm/_1060_ ;
 wire \heichips25_can_lehmann_fsm/_1061_ ;
 wire \heichips25_can_lehmann_fsm/_1062_ ;
 wire \heichips25_can_lehmann_fsm/_1063_ ;
 wire \heichips25_can_lehmann_fsm/_1064_ ;
 wire \heichips25_can_lehmann_fsm/_1065_ ;
 wire \heichips25_can_lehmann_fsm/_1066_ ;
 wire \heichips25_can_lehmann_fsm/_1067_ ;
 wire \heichips25_can_lehmann_fsm/_1068_ ;
 wire \heichips25_can_lehmann_fsm/_1069_ ;
 wire \heichips25_can_lehmann_fsm/_1070_ ;
 wire \heichips25_can_lehmann_fsm/_1071_ ;
 wire \heichips25_can_lehmann_fsm/_1072_ ;
 wire \heichips25_can_lehmann_fsm/_1073_ ;
 wire \heichips25_can_lehmann_fsm/_1074_ ;
 wire \heichips25_can_lehmann_fsm/_1075_ ;
 wire \heichips25_can_lehmann_fsm/_1076_ ;
 wire \heichips25_can_lehmann_fsm/_1077_ ;
 wire \heichips25_can_lehmann_fsm/_1078_ ;
 wire \heichips25_can_lehmann_fsm/_1079_ ;
 wire \heichips25_can_lehmann_fsm/_1080_ ;
 wire \heichips25_can_lehmann_fsm/_1081_ ;
 wire \heichips25_can_lehmann_fsm/_1082_ ;
 wire \heichips25_can_lehmann_fsm/_1083_ ;
 wire \heichips25_can_lehmann_fsm/_1084_ ;
 wire \heichips25_can_lehmann_fsm/_1085_ ;
 wire \heichips25_can_lehmann_fsm/_1086_ ;
 wire \heichips25_can_lehmann_fsm/_1087_ ;
 wire \heichips25_can_lehmann_fsm/_1088_ ;
 wire \heichips25_can_lehmann_fsm/_1089_ ;
 wire \heichips25_can_lehmann_fsm/_1090_ ;
 wire \heichips25_can_lehmann_fsm/_1091_ ;
 wire \heichips25_can_lehmann_fsm/_1092_ ;
 wire \heichips25_can_lehmann_fsm/_1093_ ;
 wire \heichips25_can_lehmann_fsm/_1094_ ;
 wire \heichips25_can_lehmann_fsm/_1095_ ;
 wire \heichips25_can_lehmann_fsm/_1096_ ;
 wire \heichips25_can_lehmann_fsm/_1097_ ;
 wire \heichips25_can_lehmann_fsm/_1098_ ;
 wire \heichips25_can_lehmann_fsm/_1099_ ;
 wire \heichips25_can_lehmann_fsm/_1100_ ;
 wire \heichips25_can_lehmann_fsm/_1101_ ;
 wire \heichips25_can_lehmann_fsm/_1102_ ;
 wire \heichips25_can_lehmann_fsm/_1103_ ;
 wire \heichips25_can_lehmann_fsm/_1104_ ;
 wire \heichips25_can_lehmann_fsm/_1105_ ;
 wire \heichips25_can_lehmann_fsm/_1106_ ;
 wire \heichips25_can_lehmann_fsm/_1107_ ;
 wire \heichips25_can_lehmann_fsm/_1108_ ;
 wire \heichips25_can_lehmann_fsm/_1109_ ;
 wire \heichips25_can_lehmann_fsm/_1110_ ;
 wire \heichips25_can_lehmann_fsm/_1111_ ;
 wire \heichips25_can_lehmann_fsm/_1112_ ;
 wire \heichips25_can_lehmann_fsm/_1113_ ;
 wire \heichips25_can_lehmann_fsm/_1114_ ;
 wire \heichips25_can_lehmann_fsm/_1115_ ;
 wire \heichips25_can_lehmann_fsm/_1116_ ;
 wire \heichips25_can_lehmann_fsm/_1117_ ;
 wire \heichips25_can_lehmann_fsm/_1118_ ;
 wire \heichips25_can_lehmann_fsm/_1119_ ;
 wire \heichips25_can_lehmann_fsm/_1120_ ;
 wire \heichips25_can_lehmann_fsm/_1121_ ;
 wire \heichips25_can_lehmann_fsm/_1122_ ;
 wire \heichips25_can_lehmann_fsm/_1123_ ;
 wire \heichips25_can_lehmann_fsm/_1124_ ;
 wire \heichips25_can_lehmann_fsm/_1125_ ;
 wire \heichips25_can_lehmann_fsm/_1126_ ;
 wire \heichips25_can_lehmann_fsm/_1127_ ;
 wire \heichips25_can_lehmann_fsm/_1128_ ;
 wire \heichips25_can_lehmann_fsm/_1129_ ;
 wire \heichips25_can_lehmann_fsm/_1130_ ;
 wire \heichips25_can_lehmann_fsm/_1131_ ;
 wire \heichips25_can_lehmann_fsm/_1132_ ;
 wire \heichips25_can_lehmann_fsm/_1133_ ;
 wire \heichips25_can_lehmann_fsm/_1134_ ;
 wire \heichips25_can_lehmann_fsm/_1135_ ;
 wire \heichips25_can_lehmann_fsm/_1136_ ;
 wire \heichips25_can_lehmann_fsm/_1137_ ;
 wire \heichips25_can_lehmann_fsm/_1138_ ;
 wire \heichips25_can_lehmann_fsm/_1139_ ;
 wire \heichips25_can_lehmann_fsm/_1140_ ;
 wire \heichips25_can_lehmann_fsm/_1141_ ;
 wire \heichips25_can_lehmann_fsm/_1142_ ;
 wire \heichips25_can_lehmann_fsm/_1143_ ;
 wire \heichips25_can_lehmann_fsm/_1144_ ;
 wire \heichips25_can_lehmann_fsm/_1145_ ;
 wire \heichips25_can_lehmann_fsm/_1146_ ;
 wire \heichips25_can_lehmann_fsm/_1147_ ;
 wire \heichips25_can_lehmann_fsm/_1148_ ;
 wire \heichips25_can_lehmann_fsm/_1149_ ;
 wire \heichips25_can_lehmann_fsm/_1150_ ;
 wire \heichips25_can_lehmann_fsm/_1151_ ;
 wire \heichips25_can_lehmann_fsm/_1152_ ;
 wire \heichips25_can_lehmann_fsm/_1153_ ;
 wire \heichips25_can_lehmann_fsm/_1154_ ;
 wire \heichips25_can_lehmann_fsm/_1155_ ;
 wire \heichips25_can_lehmann_fsm/_1156_ ;
 wire \heichips25_can_lehmann_fsm/_1157_ ;
 wire \heichips25_can_lehmann_fsm/_1158_ ;
 wire \heichips25_can_lehmann_fsm/_1159_ ;
 wire \heichips25_can_lehmann_fsm/_1160_ ;
 wire \heichips25_can_lehmann_fsm/_1161_ ;
 wire \heichips25_can_lehmann_fsm/_1162_ ;
 wire \heichips25_can_lehmann_fsm/_1163_ ;
 wire \heichips25_can_lehmann_fsm/_1164_ ;
 wire \heichips25_can_lehmann_fsm/_1165_ ;
 wire \heichips25_can_lehmann_fsm/_1166_ ;
 wire \heichips25_can_lehmann_fsm/_1167_ ;
 wire \heichips25_can_lehmann_fsm/_1168_ ;
 wire \heichips25_can_lehmann_fsm/_1169_ ;
 wire \heichips25_can_lehmann_fsm/_1170_ ;
 wire \heichips25_can_lehmann_fsm/_1171_ ;
 wire \heichips25_can_lehmann_fsm/_1172_ ;
 wire \heichips25_can_lehmann_fsm/_1173_ ;
 wire \heichips25_can_lehmann_fsm/_1174_ ;
 wire \heichips25_can_lehmann_fsm/_1175_ ;
 wire \heichips25_can_lehmann_fsm/_1176_ ;
 wire \heichips25_can_lehmann_fsm/_1177_ ;
 wire \heichips25_can_lehmann_fsm/_1178_ ;
 wire \heichips25_can_lehmann_fsm/_1179_ ;
 wire \heichips25_can_lehmann_fsm/_1180_ ;
 wire \heichips25_can_lehmann_fsm/_1181_ ;
 wire \heichips25_can_lehmann_fsm/_1182_ ;
 wire \heichips25_can_lehmann_fsm/_1183_ ;
 wire \heichips25_can_lehmann_fsm/_1184_ ;
 wire \heichips25_can_lehmann_fsm/_1185_ ;
 wire \heichips25_can_lehmann_fsm/_1186_ ;
 wire \heichips25_can_lehmann_fsm/_1187_ ;
 wire \heichips25_can_lehmann_fsm/_1188_ ;
 wire \heichips25_can_lehmann_fsm/_1189_ ;
 wire \heichips25_can_lehmann_fsm/_1190_ ;
 wire \heichips25_can_lehmann_fsm/_1191_ ;
 wire \heichips25_can_lehmann_fsm/_1192_ ;
 wire \heichips25_can_lehmann_fsm/_1193_ ;
 wire \heichips25_can_lehmann_fsm/_1194_ ;
 wire \heichips25_can_lehmann_fsm/_1195_ ;
 wire \heichips25_can_lehmann_fsm/_1196_ ;
 wire \heichips25_can_lehmann_fsm/_1197_ ;
 wire \heichips25_can_lehmann_fsm/_1198_ ;
 wire \heichips25_can_lehmann_fsm/_1199_ ;
 wire \heichips25_can_lehmann_fsm/_1200_ ;
 wire \heichips25_can_lehmann_fsm/_1201_ ;
 wire \heichips25_can_lehmann_fsm/_1202_ ;
 wire \heichips25_can_lehmann_fsm/_1203_ ;
 wire \heichips25_can_lehmann_fsm/_1204_ ;
 wire \heichips25_can_lehmann_fsm/_1205_ ;
 wire \heichips25_can_lehmann_fsm/_1206_ ;
 wire \heichips25_can_lehmann_fsm/_1207_ ;
 wire \heichips25_can_lehmann_fsm/_1208_ ;
 wire \heichips25_can_lehmann_fsm/_1209_ ;
 wire \heichips25_can_lehmann_fsm/_1210_ ;
 wire \heichips25_can_lehmann_fsm/_1211_ ;
 wire \heichips25_can_lehmann_fsm/_1212_ ;
 wire \heichips25_can_lehmann_fsm/_1213_ ;
 wire \heichips25_can_lehmann_fsm/_1214_ ;
 wire \heichips25_can_lehmann_fsm/_1215_ ;
 wire \heichips25_can_lehmann_fsm/_1216_ ;
 wire \heichips25_can_lehmann_fsm/_1217_ ;
 wire \heichips25_can_lehmann_fsm/_1218_ ;
 wire \heichips25_can_lehmann_fsm/_1219_ ;
 wire \heichips25_can_lehmann_fsm/_1220_ ;
 wire \heichips25_can_lehmann_fsm/_1221_ ;
 wire \heichips25_can_lehmann_fsm/_1222_ ;
 wire \heichips25_can_lehmann_fsm/_1223_ ;
 wire \heichips25_can_lehmann_fsm/_1224_ ;
 wire \heichips25_can_lehmann_fsm/_1225_ ;
 wire \heichips25_can_lehmann_fsm/_1226_ ;
 wire \heichips25_can_lehmann_fsm/_1227_ ;
 wire \heichips25_can_lehmann_fsm/_1228_ ;
 wire \heichips25_can_lehmann_fsm/_1229_ ;
 wire \heichips25_can_lehmann_fsm/_1230_ ;
 wire \heichips25_can_lehmann_fsm/_1231_ ;
 wire \heichips25_can_lehmann_fsm/_1232_ ;
 wire \heichips25_can_lehmann_fsm/_1233_ ;
 wire \heichips25_can_lehmann_fsm/_1234_ ;
 wire \heichips25_can_lehmann_fsm/_1235_ ;
 wire \heichips25_can_lehmann_fsm/_1236_ ;
 wire \heichips25_can_lehmann_fsm/_1237_ ;
 wire \heichips25_can_lehmann_fsm/_1238_ ;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire \heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[0] ;
 wire \heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[10] ;
 wire \heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[11] ;
 wire \heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[12] ;
 wire \heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[13] ;
 wire \heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[14] ;
 wire \heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[15] ;
 wire \heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[16] ;
 wire \heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[17] ;
 wire \heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[18] ;
 wire \heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[19] ;
 wire \heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[1] ;
 wire \heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[20] ;
 wire \heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[21] ;
 wire \heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[22] ;
 wire \heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[23] ;
 wire \heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[2] ;
 wire \heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[3] ;
 wire \heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[4] ;
 wire \heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[5] ;
 wire \heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[6] ;
 wire \heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[7] ;
 wire \heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[8] ;
 wire \heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[9] ;
 wire \heichips25_can_lehmann_fsm/controller.const_data[0] ;
 wire \heichips25_can_lehmann_fsm/controller.const_data[10] ;
 wire \heichips25_can_lehmann_fsm/controller.const_data[11] ;
 wire \heichips25_can_lehmann_fsm/controller.const_data[12] ;
 wire \heichips25_can_lehmann_fsm/controller.const_data[13] ;
 wire \heichips25_can_lehmann_fsm/controller.const_data[14] ;
 wire \heichips25_can_lehmann_fsm/controller.const_data[15] ;
 wire \heichips25_can_lehmann_fsm/controller.const_data[16] ;
 wire \heichips25_can_lehmann_fsm/controller.const_data[17] ;
 wire \heichips25_can_lehmann_fsm/controller.const_data[18] ;
 wire \heichips25_can_lehmann_fsm/controller.const_data[19] ;
 wire \heichips25_can_lehmann_fsm/controller.const_data[1] ;
 wire \heichips25_can_lehmann_fsm/controller.const_data[20] ;
 wire \heichips25_can_lehmann_fsm/controller.const_data[21] ;
 wire \heichips25_can_lehmann_fsm/controller.const_data[22] ;
 wire \heichips25_can_lehmann_fsm/controller.const_data[23] ;
 wire \heichips25_can_lehmann_fsm/controller.const_data[24] ;
 wire \heichips25_can_lehmann_fsm/controller.const_data[25] ;
 wire \heichips25_can_lehmann_fsm/controller.const_data[26] ;
 wire \heichips25_can_lehmann_fsm/controller.const_data[27] ;
 wire \heichips25_can_lehmann_fsm/controller.const_data[28] ;
 wire \heichips25_can_lehmann_fsm/controller.const_data[29] ;
 wire \heichips25_can_lehmann_fsm/controller.const_data[2] ;
 wire \heichips25_can_lehmann_fsm/controller.const_data[30] ;
 wire \heichips25_can_lehmann_fsm/controller.const_data[31] ;
 wire \heichips25_can_lehmann_fsm/controller.const_data[3] ;
 wire \heichips25_can_lehmann_fsm/controller.const_data[4] ;
 wire \heichips25_can_lehmann_fsm/controller.const_data[5] ;
 wire \heichips25_can_lehmann_fsm/controller.const_data[6] ;
 wire \heichips25_can_lehmann_fsm/controller.const_data[7] ;
 wire \heichips25_can_lehmann_fsm/controller.const_data[8] ;
 wire \heichips25_can_lehmann_fsm/controller.const_data[9] ;
 wire \heichips25_can_lehmann_fsm/controller.counter2.counter_0[0] ;
 wire \heichips25_can_lehmann_fsm/controller.counter2.counter_0[10] ;
 wire \heichips25_can_lehmann_fsm/controller.counter2.counter_0[11] ;
 wire \heichips25_can_lehmann_fsm/controller.counter2.counter_0[12] ;
 wire \heichips25_can_lehmann_fsm/controller.counter2.counter_0[13] ;
 wire \heichips25_can_lehmann_fsm/controller.counter2.counter_0[14] ;
 wire \heichips25_can_lehmann_fsm/controller.counter2.counter_0[15] ;
 wire \heichips25_can_lehmann_fsm/controller.counter2.counter_0[1] ;
 wire \heichips25_can_lehmann_fsm/controller.counter2.counter_0[2] ;
 wire \heichips25_can_lehmann_fsm/controller.counter2.counter_0[3] ;
 wire \heichips25_can_lehmann_fsm/controller.counter2.counter_0[4] ;
 wire \heichips25_can_lehmann_fsm/controller.counter2.counter_0[5] ;
 wire \heichips25_can_lehmann_fsm/controller.counter2.counter_0[6] ;
 wire \heichips25_can_lehmann_fsm/controller.counter2.counter_0[7] ;
 wire \heichips25_can_lehmann_fsm/controller.counter2.counter_0[8] ;
 wire \heichips25_can_lehmann_fsm/controller.counter2.counter_0[9] ;
 wire \heichips25_can_lehmann_fsm/controller.counter2.counter_1[0] ;
 wire \heichips25_can_lehmann_fsm/controller.counter2.counter_1[10] ;
 wire \heichips25_can_lehmann_fsm/controller.counter2.counter_1[11] ;
 wire \heichips25_can_lehmann_fsm/controller.counter2.counter_1[12] ;
 wire \heichips25_can_lehmann_fsm/controller.counter2.counter_1[13] ;
 wire \heichips25_can_lehmann_fsm/controller.counter2.counter_1[14] ;
 wire \heichips25_can_lehmann_fsm/controller.counter2.counter_1[15] ;
 wire \heichips25_can_lehmann_fsm/controller.counter2.counter_1[1] ;
 wire \heichips25_can_lehmann_fsm/controller.counter2.counter_1[2] ;
 wire \heichips25_can_lehmann_fsm/controller.counter2.counter_1[3] ;
 wire \heichips25_can_lehmann_fsm/controller.counter2.counter_1[4] ;
 wire \heichips25_can_lehmann_fsm/controller.counter2.counter_1[5] ;
 wire \heichips25_can_lehmann_fsm/controller.counter2.counter_1[6] ;
 wire \heichips25_can_lehmann_fsm/controller.counter2.counter_1[7] ;
 wire \heichips25_can_lehmann_fsm/controller.counter2.counter_1[8] ;
 wire \heichips25_can_lehmann_fsm/controller.counter2.counter_1[9] ;
 wire \heichips25_can_lehmann_fsm/controller.extended_cond.opcode[0] ;
 wire \heichips25_can_lehmann_fsm/controller.extended_cond.opcode[1] ;
 wire \heichips25_can_lehmann_fsm/controller.extended_cond.opcode[2] ;
 wire \heichips25_can_lehmann_fsm/controller.extended_jump_target[0] ;
 wire \heichips25_can_lehmann_fsm/controller.extended_jump_target[1] ;
 wire \heichips25_can_lehmann_fsm/controller.extended_jump_target[2] ;
 wire \heichips25_can_lehmann_fsm/controller.extended_state[0] ;
 wire \heichips25_can_lehmann_fsm/controller.extended_state[1] ;
 wire \heichips25_can_lehmann_fsm/controller.extended_state[2] ;
 wire \heichips25_can_lehmann_fsm/controller.extended_then_action[0] ;
 wire \heichips25_can_lehmann_fsm/controller.extended_then_action[1] ;
 wire \heichips25_can_lehmann_fsm/controller.extended_then_action[2] ;
 wire \heichips25_can_lehmann_fsm/controller.extended_then_action[3] ;
 wire \heichips25_can_lehmann_fsm/controller.extended_then_action[4] ;
 wire \heichips25_can_lehmann_fsm/controller.extended_then_action[5] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.addr[0] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.addr[1] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.addr[2] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[18] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[19] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[20] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[21] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[22] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[23] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[3] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[4] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[5] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[6] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[7] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[8] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[100] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[101] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[102] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[103] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[104] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[105] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[106] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[107] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[108] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[109] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[110] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[111] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[112] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[113] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[114] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[115] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[116] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[117] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[118] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[119] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[120] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[121] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[122] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[123] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[124] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[125] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[126] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[127] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[128] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[129] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[130] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[131] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[132] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[133] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[134] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[135] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[136] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[137] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[138] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[139] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[140] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[141] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[142] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[143] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[144] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[145] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[146] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[147] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[148] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[149] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[150] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[151] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[152] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[153] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[154] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[155] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[156] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[157] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[158] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[159] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[160] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[161] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[162] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[163] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[164] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[165] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[166] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[167] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[168] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[169] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[170] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[171] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[172] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[173] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[174] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[175] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[176] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[177] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[178] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[179] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[180] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[181] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[182] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[183] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[184] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[185] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[186] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[187] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[188] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[189] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[190] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[191] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[192] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[193] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[194] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[195] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[196] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[197] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[198] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[199] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[32] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[33] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[34] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[35] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[36] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[37] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[38] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[39] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[40] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[41] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[42] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[43] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[44] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[45] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[46] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[47] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[48] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[49] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[50] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[51] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[52] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[53] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[54] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[55] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[56] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[57] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[58] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[59] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[60] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[61] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[62] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[63] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[64] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[65] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[66] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[67] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[68] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[69] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[70] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[71] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[72] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[73] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[74] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[75] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[76] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[77] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[78] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[79] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[80] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[81] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[82] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[83] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[84] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[85] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[86] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[87] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[88] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[89] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[90] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[91] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[92] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[93] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[94] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[95] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[96] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[97] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[98] ;
 wire \heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[99] ;
 wire \heichips25_can_lehmann_fsm/controller.output_controller.keep[0] ;
 wire \heichips25_can_lehmann_fsm/controller.output_controller.keep[1] ;
 wire \heichips25_can_lehmann_fsm/controller.output_controller.keep[2] ;
 wire \heichips25_sap3/_0000_ ;
 wire \heichips25_sap3/_0001_ ;
 wire \heichips25_sap3/_0002_ ;
 wire \heichips25_sap3/_0003_ ;
 wire \heichips25_sap3/_0004_ ;
 wire \heichips25_sap3/_0005_ ;
 wire \heichips25_sap3/_0006_ ;
 wire \heichips25_sap3/_0007_ ;
 wire \heichips25_sap3/_0008_ ;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire \heichips25_sap3/_0017_ ;
 wire \heichips25_sap3/_0018_ ;
 wire net823;
 wire net824;
 wire net825;
 wire clknet_leaf_0_clk;
 wire \heichips25_sap3/_0023_ ;
 wire \heichips25_sap3/_0024_ ;
 wire \heichips25_sap3/_0025_ ;
 wire \heichips25_sap3/_0026_ ;
 wire \heichips25_sap3/_0027_ ;
 wire \heichips25_sap3/_0028_ ;
 wire \heichips25_sap3/_0029_ ;
 wire \heichips25_sap3/_0030_ ;
 wire \heichips25_sap3/_0031_ ;
 wire \heichips25_sap3/_0032_ ;
 wire \heichips25_sap3/_0033_ ;
 wire \heichips25_sap3/_0034_ ;
 wire \heichips25_sap3/_0035_ ;
 wire \heichips25_sap3/_0036_ ;
 wire \heichips25_sap3/_0037_ ;
 wire \heichips25_sap3/_0038_ ;
 wire \heichips25_sap3/_0039_ ;
 wire \heichips25_sap3/_0040_ ;
 wire \heichips25_sap3/_0041_ ;
 wire \heichips25_sap3/_0042_ ;
 wire \heichips25_sap3/_0043_ ;
 wire \heichips25_sap3/_0044_ ;
 wire \heichips25_sap3/_0045_ ;
 wire \heichips25_sap3/_0046_ ;
 wire \heichips25_sap3/_0047_ ;
 wire \heichips25_sap3/_0048_ ;
 wire \heichips25_sap3/_0049_ ;
 wire \heichips25_sap3/_0050_ ;
 wire \heichips25_sap3/_0051_ ;
 wire \heichips25_sap3/_0052_ ;
 wire \heichips25_sap3/_0053_ ;
 wire \heichips25_sap3/_0054_ ;
 wire \heichips25_sap3/_0055_ ;
 wire \heichips25_sap3/_0056_ ;
 wire \heichips25_sap3/_0057_ ;
 wire \heichips25_sap3/_0058_ ;
 wire \heichips25_sap3/_0059_ ;
 wire \heichips25_sap3/_0060_ ;
 wire \heichips25_sap3/_0061_ ;
 wire \heichips25_sap3/_0062_ ;
 wire \heichips25_sap3/_0063_ ;
 wire \heichips25_sap3/_0064_ ;
 wire \heichips25_sap3/_0065_ ;
 wire \heichips25_sap3/_0066_ ;
 wire \heichips25_sap3/_0067_ ;
 wire \heichips25_sap3/_0068_ ;
 wire \heichips25_sap3/_0069_ ;
 wire \heichips25_sap3/_0070_ ;
 wire \heichips25_sap3/_0071_ ;
 wire \heichips25_sap3/_0072_ ;
 wire \heichips25_sap3/_0073_ ;
 wire \heichips25_sap3/_0074_ ;
 wire \heichips25_sap3/_0075_ ;
 wire \heichips25_sap3/_0076_ ;
 wire \heichips25_sap3/_0077_ ;
 wire \heichips25_sap3/_0078_ ;
 wire \heichips25_sap3/_0079_ ;
 wire \heichips25_sap3/_0080_ ;
 wire \heichips25_sap3/_0081_ ;
 wire \heichips25_sap3/_0082_ ;
 wire \heichips25_sap3/_0083_ ;
 wire \heichips25_sap3/_0084_ ;
 wire \heichips25_sap3/_0085_ ;
 wire \heichips25_sap3/_0086_ ;
 wire \heichips25_sap3/_0087_ ;
 wire \heichips25_sap3/_0088_ ;
 wire \heichips25_sap3/_0089_ ;
 wire \heichips25_sap3/_0090_ ;
 wire \heichips25_sap3/_0091_ ;
 wire \heichips25_sap3/_0092_ ;
 wire \heichips25_sap3/_0093_ ;
 wire \heichips25_sap3/_0094_ ;
 wire \heichips25_sap3/_0095_ ;
 wire \heichips25_sap3/_0096_ ;
 wire \heichips25_sap3/_0097_ ;
 wire \heichips25_sap3/_0098_ ;
 wire \heichips25_sap3/_0099_ ;
 wire \heichips25_sap3/_0100_ ;
 wire \heichips25_sap3/_0101_ ;
 wire \heichips25_sap3/_0102_ ;
 wire \heichips25_sap3/_0103_ ;
 wire \heichips25_sap3/_0104_ ;
 wire \heichips25_sap3/_0105_ ;
 wire \heichips25_sap3/_0106_ ;
 wire \heichips25_sap3/_0107_ ;
 wire \heichips25_sap3/_0108_ ;
 wire \heichips25_sap3/_0109_ ;
 wire \heichips25_sap3/_0110_ ;
 wire \heichips25_sap3/_0111_ ;
 wire \heichips25_sap3/_0112_ ;
 wire \heichips25_sap3/_0113_ ;
 wire \heichips25_sap3/_0114_ ;
 wire \heichips25_sap3/_0115_ ;
 wire \heichips25_sap3/_0116_ ;
 wire \heichips25_sap3/_0117_ ;
 wire \heichips25_sap3/_0118_ ;
 wire \heichips25_sap3/_0119_ ;
 wire \heichips25_sap3/_0120_ ;
 wire \heichips25_sap3/_0121_ ;
 wire \heichips25_sap3/_0122_ ;
 wire \heichips25_sap3/_0123_ ;
 wire \heichips25_sap3/_0124_ ;
 wire \heichips25_sap3/_0125_ ;
 wire \heichips25_sap3/_0126_ ;
 wire \heichips25_sap3/_0127_ ;
 wire \heichips25_sap3/_0128_ ;
 wire \heichips25_sap3/_0129_ ;
 wire \heichips25_sap3/_0130_ ;
 wire \heichips25_sap3/_0131_ ;
 wire \heichips25_sap3/_0132_ ;
 wire \heichips25_sap3/_0133_ ;
 wire \heichips25_sap3/_0134_ ;
 wire \heichips25_sap3/_0135_ ;
 wire \heichips25_sap3/_0136_ ;
 wire \heichips25_sap3/_0137_ ;
 wire \heichips25_sap3/_0138_ ;
 wire \heichips25_sap3/_0139_ ;
 wire \heichips25_sap3/_0140_ ;
 wire \heichips25_sap3/_0141_ ;
 wire \heichips25_sap3/_0142_ ;
 wire \heichips25_sap3/_0143_ ;
 wire \heichips25_sap3/_0144_ ;
 wire \heichips25_sap3/_0145_ ;
 wire \heichips25_sap3/_0146_ ;
 wire \heichips25_sap3/_0147_ ;
 wire \heichips25_sap3/_0148_ ;
 wire \heichips25_sap3/_0149_ ;
 wire \heichips25_sap3/_0150_ ;
 wire \heichips25_sap3/_0151_ ;
 wire \heichips25_sap3/_0152_ ;
 wire \heichips25_sap3/_0153_ ;
 wire \heichips25_sap3/_0154_ ;
 wire \heichips25_sap3/_0155_ ;
 wire \heichips25_sap3/_0156_ ;
 wire \heichips25_sap3/_0157_ ;
 wire \heichips25_sap3/_0158_ ;
 wire \heichips25_sap3/_0159_ ;
 wire \heichips25_sap3/_0160_ ;
 wire \heichips25_sap3/_0161_ ;
 wire \heichips25_sap3/_0162_ ;
 wire \heichips25_sap3/_0163_ ;
 wire \heichips25_sap3/_0164_ ;
 wire \heichips25_sap3/_0165_ ;
 wire \heichips25_sap3/_0166_ ;
 wire \heichips25_sap3/_0167_ ;
 wire \heichips25_sap3/_0168_ ;
 wire \heichips25_sap3/_0169_ ;
 wire \heichips25_sap3/_0170_ ;
 wire \heichips25_sap3/_0171_ ;
 wire \heichips25_sap3/_0172_ ;
 wire \heichips25_sap3/_0173_ ;
 wire \heichips25_sap3/_0174_ ;
 wire \heichips25_sap3/_0175_ ;
 wire \heichips25_sap3/_0176_ ;
 wire \heichips25_sap3/_0177_ ;
 wire \heichips25_sap3/_0178_ ;
 wire \heichips25_sap3/_0179_ ;
 wire \heichips25_sap3/_0180_ ;
 wire \heichips25_sap3/_0181_ ;
 wire \heichips25_sap3/_0182_ ;
 wire \heichips25_sap3/_0183_ ;
 wire \heichips25_sap3/_0184_ ;
 wire \heichips25_sap3/_0185_ ;
 wire \heichips25_sap3/_0186_ ;
 wire \heichips25_sap3/_0187_ ;
 wire \heichips25_sap3/_0188_ ;
 wire \heichips25_sap3/_0189_ ;
 wire \heichips25_sap3/_0190_ ;
 wire \heichips25_sap3/_0191_ ;
 wire \heichips25_sap3/_0192_ ;
 wire \heichips25_sap3/_0193_ ;
 wire \heichips25_sap3/_0194_ ;
 wire \heichips25_sap3/_0195_ ;
 wire \heichips25_sap3/_0196_ ;
 wire \heichips25_sap3/_0197_ ;
 wire \heichips25_sap3/_0198_ ;
 wire \heichips25_sap3/_0199_ ;
 wire \heichips25_sap3/_0200_ ;
 wire \heichips25_sap3/_0201_ ;
 wire \heichips25_sap3/_0202_ ;
 wire \heichips25_sap3/_0203_ ;
 wire \heichips25_sap3/_0204_ ;
 wire \heichips25_sap3/_0205_ ;
 wire \heichips25_sap3/_0206_ ;
 wire \heichips25_sap3/_0207_ ;
 wire \heichips25_sap3/_0208_ ;
 wire \heichips25_sap3/_0209_ ;
 wire \heichips25_sap3/_0210_ ;
 wire \heichips25_sap3/_0211_ ;
 wire \heichips25_sap3/_0212_ ;
 wire \heichips25_sap3/_0213_ ;
 wire \heichips25_sap3/_0214_ ;
 wire \heichips25_sap3/_0215_ ;
 wire \heichips25_sap3/_0216_ ;
 wire \heichips25_sap3/_0217_ ;
 wire \heichips25_sap3/_0218_ ;
 wire \heichips25_sap3/_0219_ ;
 wire \heichips25_sap3/_0220_ ;
 wire \heichips25_sap3/_0221_ ;
 wire \heichips25_sap3/_0222_ ;
 wire \heichips25_sap3/_0223_ ;
 wire \heichips25_sap3/_0224_ ;
 wire \heichips25_sap3/_0225_ ;
 wire \heichips25_sap3/_0226_ ;
 wire \heichips25_sap3/_0227_ ;
 wire \heichips25_sap3/_0228_ ;
 wire \heichips25_sap3/_0229_ ;
 wire \heichips25_sap3/_0230_ ;
 wire \heichips25_sap3/_0231_ ;
 wire \heichips25_sap3/_0232_ ;
 wire \heichips25_sap3/_0233_ ;
 wire \heichips25_sap3/_0234_ ;
 wire \heichips25_sap3/_0235_ ;
 wire \heichips25_sap3/_0236_ ;
 wire \heichips25_sap3/_0237_ ;
 wire \heichips25_sap3/_0238_ ;
 wire \heichips25_sap3/_0239_ ;
 wire \heichips25_sap3/_0240_ ;
 wire \heichips25_sap3/_0241_ ;
 wire \heichips25_sap3/_0242_ ;
 wire \heichips25_sap3/_0243_ ;
 wire \heichips25_sap3/_0244_ ;
 wire \heichips25_sap3/_0245_ ;
 wire \heichips25_sap3/_0246_ ;
 wire \heichips25_sap3/_0247_ ;
 wire \heichips25_sap3/_0248_ ;
 wire \heichips25_sap3/_0249_ ;
 wire \heichips25_sap3/_0250_ ;
 wire \heichips25_sap3/_0251_ ;
 wire \heichips25_sap3/_0252_ ;
 wire \heichips25_sap3/_0253_ ;
 wire \heichips25_sap3/_0254_ ;
 wire \heichips25_sap3/_0255_ ;
 wire \heichips25_sap3/_0256_ ;
 wire \heichips25_sap3/_0257_ ;
 wire \heichips25_sap3/_0258_ ;
 wire \heichips25_sap3/_0259_ ;
 wire \heichips25_sap3/_0260_ ;
 wire \heichips25_sap3/_0261_ ;
 wire \heichips25_sap3/_0262_ ;
 wire \heichips25_sap3/_0263_ ;
 wire \heichips25_sap3/_0264_ ;
 wire \heichips25_sap3/_0265_ ;
 wire \heichips25_sap3/_0266_ ;
 wire \heichips25_sap3/_0267_ ;
 wire \heichips25_sap3/_0268_ ;
 wire \heichips25_sap3/_0269_ ;
 wire \heichips25_sap3/_0270_ ;
 wire \heichips25_sap3/_0271_ ;
 wire \heichips25_sap3/_0272_ ;
 wire \heichips25_sap3/_0273_ ;
 wire \heichips25_sap3/_0274_ ;
 wire \heichips25_sap3/_0275_ ;
 wire \heichips25_sap3/_0276_ ;
 wire \heichips25_sap3/_0277_ ;
 wire \heichips25_sap3/_0278_ ;
 wire \heichips25_sap3/_0279_ ;
 wire \heichips25_sap3/_0280_ ;
 wire \heichips25_sap3/_0281_ ;
 wire \heichips25_sap3/_0282_ ;
 wire \heichips25_sap3/_0283_ ;
 wire \heichips25_sap3/_0284_ ;
 wire \heichips25_sap3/_0285_ ;
 wire \heichips25_sap3/_0286_ ;
 wire \heichips25_sap3/_0287_ ;
 wire \heichips25_sap3/_0288_ ;
 wire \heichips25_sap3/_0289_ ;
 wire \heichips25_sap3/_0290_ ;
 wire \heichips25_sap3/_0291_ ;
 wire \heichips25_sap3/_0292_ ;
 wire \heichips25_sap3/_0293_ ;
 wire \heichips25_sap3/_0294_ ;
 wire \heichips25_sap3/_0295_ ;
 wire \heichips25_sap3/_0296_ ;
 wire \heichips25_sap3/_0297_ ;
 wire \heichips25_sap3/_0298_ ;
 wire \heichips25_sap3/_0299_ ;
 wire \heichips25_sap3/_0300_ ;
 wire \heichips25_sap3/_0301_ ;
 wire \heichips25_sap3/_0302_ ;
 wire \heichips25_sap3/_0303_ ;
 wire \heichips25_sap3/_0304_ ;
 wire \heichips25_sap3/_0305_ ;
 wire \heichips25_sap3/_0306_ ;
 wire \heichips25_sap3/_0307_ ;
 wire \heichips25_sap3/_0308_ ;
 wire \heichips25_sap3/_0309_ ;
 wire \heichips25_sap3/_0310_ ;
 wire \heichips25_sap3/_0311_ ;
 wire \heichips25_sap3/_0312_ ;
 wire \heichips25_sap3/_0313_ ;
 wire \heichips25_sap3/_0314_ ;
 wire \heichips25_sap3/_0315_ ;
 wire \heichips25_sap3/_0316_ ;
 wire \heichips25_sap3/_0317_ ;
 wire \heichips25_sap3/_0318_ ;
 wire \heichips25_sap3/_0319_ ;
 wire \heichips25_sap3/_0320_ ;
 wire \heichips25_sap3/_0321_ ;
 wire \heichips25_sap3/_0322_ ;
 wire \heichips25_sap3/_0323_ ;
 wire \heichips25_sap3/_0324_ ;
 wire \heichips25_sap3/_0325_ ;
 wire \heichips25_sap3/_0326_ ;
 wire \heichips25_sap3/_0327_ ;
 wire \heichips25_sap3/_0328_ ;
 wire \heichips25_sap3/_0329_ ;
 wire \heichips25_sap3/_0330_ ;
 wire \heichips25_sap3/_0331_ ;
 wire \heichips25_sap3/_0332_ ;
 wire \heichips25_sap3/_0333_ ;
 wire \heichips25_sap3/_0334_ ;
 wire \heichips25_sap3/_0335_ ;
 wire \heichips25_sap3/_0336_ ;
 wire \heichips25_sap3/_0337_ ;
 wire \heichips25_sap3/_0338_ ;
 wire \heichips25_sap3/_0339_ ;
 wire \heichips25_sap3/_0340_ ;
 wire \heichips25_sap3/_0341_ ;
 wire \heichips25_sap3/_0342_ ;
 wire \heichips25_sap3/_0343_ ;
 wire \heichips25_sap3/_0344_ ;
 wire \heichips25_sap3/_0345_ ;
 wire \heichips25_sap3/_0346_ ;
 wire \heichips25_sap3/_0347_ ;
 wire \heichips25_sap3/_0348_ ;
 wire \heichips25_sap3/_0349_ ;
 wire \heichips25_sap3/_0350_ ;
 wire \heichips25_sap3/_0351_ ;
 wire \heichips25_sap3/_0352_ ;
 wire \heichips25_sap3/_0353_ ;
 wire \heichips25_sap3/_0354_ ;
 wire \heichips25_sap3/_0355_ ;
 wire \heichips25_sap3/_0356_ ;
 wire \heichips25_sap3/_0357_ ;
 wire \heichips25_sap3/_0358_ ;
 wire \heichips25_sap3/_0359_ ;
 wire \heichips25_sap3/_0360_ ;
 wire \heichips25_sap3/_0361_ ;
 wire \heichips25_sap3/_0362_ ;
 wire \heichips25_sap3/_0363_ ;
 wire \heichips25_sap3/_0364_ ;
 wire \heichips25_sap3/_0365_ ;
 wire \heichips25_sap3/_0366_ ;
 wire \heichips25_sap3/_0367_ ;
 wire \heichips25_sap3/_0368_ ;
 wire \heichips25_sap3/_0369_ ;
 wire \heichips25_sap3/_0370_ ;
 wire \heichips25_sap3/_0371_ ;
 wire \heichips25_sap3/_0372_ ;
 wire \heichips25_sap3/_0373_ ;
 wire \heichips25_sap3/_0374_ ;
 wire \heichips25_sap3/_0375_ ;
 wire \heichips25_sap3/_0376_ ;
 wire \heichips25_sap3/_0377_ ;
 wire \heichips25_sap3/_0378_ ;
 wire \heichips25_sap3/_0379_ ;
 wire \heichips25_sap3/_0380_ ;
 wire \heichips25_sap3/_0381_ ;
 wire \heichips25_sap3/_0382_ ;
 wire \heichips25_sap3/_0383_ ;
 wire \heichips25_sap3/_0384_ ;
 wire \heichips25_sap3/_0385_ ;
 wire \heichips25_sap3/_0386_ ;
 wire \heichips25_sap3/_0387_ ;
 wire \heichips25_sap3/_0388_ ;
 wire \heichips25_sap3/_0389_ ;
 wire \heichips25_sap3/_0390_ ;
 wire \heichips25_sap3/_0391_ ;
 wire \heichips25_sap3/_0392_ ;
 wire \heichips25_sap3/_0393_ ;
 wire \heichips25_sap3/_0394_ ;
 wire \heichips25_sap3/_0395_ ;
 wire \heichips25_sap3/_0396_ ;
 wire \heichips25_sap3/_0397_ ;
 wire \heichips25_sap3/_0398_ ;
 wire \heichips25_sap3/_0399_ ;
 wire \heichips25_sap3/_0400_ ;
 wire \heichips25_sap3/_0401_ ;
 wire \heichips25_sap3/_0402_ ;
 wire \heichips25_sap3/_0403_ ;
 wire \heichips25_sap3/_0404_ ;
 wire \heichips25_sap3/_0405_ ;
 wire \heichips25_sap3/_0406_ ;
 wire \heichips25_sap3/_0407_ ;
 wire \heichips25_sap3/_0408_ ;
 wire \heichips25_sap3/_0409_ ;
 wire \heichips25_sap3/_0410_ ;
 wire \heichips25_sap3/_0411_ ;
 wire \heichips25_sap3/_0412_ ;
 wire \heichips25_sap3/_0413_ ;
 wire \heichips25_sap3/_0414_ ;
 wire \heichips25_sap3/_0415_ ;
 wire \heichips25_sap3/_0416_ ;
 wire \heichips25_sap3/_0417_ ;
 wire \heichips25_sap3/_0418_ ;
 wire \heichips25_sap3/_0419_ ;
 wire \heichips25_sap3/_0420_ ;
 wire \heichips25_sap3/_0421_ ;
 wire \heichips25_sap3/_0422_ ;
 wire \heichips25_sap3/_0423_ ;
 wire \heichips25_sap3/_0424_ ;
 wire \heichips25_sap3/_0425_ ;
 wire \heichips25_sap3/_0426_ ;
 wire \heichips25_sap3/_0427_ ;
 wire \heichips25_sap3/_0428_ ;
 wire \heichips25_sap3/_0429_ ;
 wire \heichips25_sap3/_0430_ ;
 wire \heichips25_sap3/_0431_ ;
 wire \heichips25_sap3/_0432_ ;
 wire \heichips25_sap3/_0433_ ;
 wire \heichips25_sap3/_0434_ ;
 wire \heichips25_sap3/_0435_ ;
 wire \heichips25_sap3/_0436_ ;
 wire \heichips25_sap3/_0437_ ;
 wire \heichips25_sap3/_0438_ ;
 wire \heichips25_sap3/_0439_ ;
 wire \heichips25_sap3/_0440_ ;
 wire \heichips25_sap3/_0441_ ;
 wire \heichips25_sap3/_0442_ ;
 wire \heichips25_sap3/_0443_ ;
 wire \heichips25_sap3/_0444_ ;
 wire \heichips25_sap3/_0445_ ;
 wire \heichips25_sap3/_0446_ ;
 wire \heichips25_sap3/_0447_ ;
 wire \heichips25_sap3/_0448_ ;
 wire \heichips25_sap3/_0449_ ;
 wire \heichips25_sap3/_0450_ ;
 wire \heichips25_sap3/_0451_ ;
 wire \heichips25_sap3/_0452_ ;
 wire \heichips25_sap3/_0453_ ;
 wire \heichips25_sap3/_0454_ ;
 wire \heichips25_sap3/_0455_ ;
 wire \heichips25_sap3/_0456_ ;
 wire \heichips25_sap3/_0457_ ;
 wire \heichips25_sap3/_0458_ ;
 wire \heichips25_sap3/_0459_ ;
 wire \heichips25_sap3/_0460_ ;
 wire \heichips25_sap3/_0461_ ;
 wire \heichips25_sap3/_0462_ ;
 wire \heichips25_sap3/_0463_ ;
 wire \heichips25_sap3/_0464_ ;
 wire \heichips25_sap3/_0465_ ;
 wire \heichips25_sap3/_0466_ ;
 wire \heichips25_sap3/_0467_ ;
 wire \heichips25_sap3/_0468_ ;
 wire \heichips25_sap3/_0469_ ;
 wire \heichips25_sap3/_0470_ ;
 wire \heichips25_sap3/_0471_ ;
 wire \heichips25_sap3/_0472_ ;
 wire \heichips25_sap3/_0473_ ;
 wire \heichips25_sap3/_0474_ ;
 wire \heichips25_sap3/_0475_ ;
 wire \heichips25_sap3/_0476_ ;
 wire \heichips25_sap3/_0477_ ;
 wire \heichips25_sap3/_0478_ ;
 wire \heichips25_sap3/_0479_ ;
 wire \heichips25_sap3/_0480_ ;
 wire \heichips25_sap3/_0481_ ;
 wire \heichips25_sap3/_0482_ ;
 wire \heichips25_sap3/_0483_ ;
 wire \heichips25_sap3/_0484_ ;
 wire \heichips25_sap3/_0485_ ;
 wire \heichips25_sap3/_0486_ ;
 wire \heichips25_sap3/_0487_ ;
 wire \heichips25_sap3/_0488_ ;
 wire \heichips25_sap3/_0489_ ;
 wire \heichips25_sap3/_0490_ ;
 wire \heichips25_sap3/_0491_ ;
 wire \heichips25_sap3/_0492_ ;
 wire \heichips25_sap3/_0493_ ;
 wire \heichips25_sap3/_0494_ ;
 wire \heichips25_sap3/_0495_ ;
 wire \heichips25_sap3/_0496_ ;
 wire \heichips25_sap3/_0497_ ;
 wire \heichips25_sap3/_0498_ ;
 wire \heichips25_sap3/_0499_ ;
 wire \heichips25_sap3/_0500_ ;
 wire \heichips25_sap3/_0501_ ;
 wire \heichips25_sap3/_0502_ ;
 wire \heichips25_sap3/_0503_ ;
 wire \heichips25_sap3/_0504_ ;
 wire \heichips25_sap3/_0505_ ;
 wire \heichips25_sap3/_0506_ ;
 wire \heichips25_sap3/_0507_ ;
 wire \heichips25_sap3/_0508_ ;
 wire \heichips25_sap3/_0509_ ;
 wire \heichips25_sap3/_0510_ ;
 wire \heichips25_sap3/_0511_ ;
 wire \heichips25_sap3/_0512_ ;
 wire \heichips25_sap3/_0513_ ;
 wire \heichips25_sap3/_0514_ ;
 wire \heichips25_sap3/_0515_ ;
 wire \heichips25_sap3/_0516_ ;
 wire \heichips25_sap3/_0517_ ;
 wire \heichips25_sap3/_0518_ ;
 wire \heichips25_sap3/_0519_ ;
 wire \heichips25_sap3/_0520_ ;
 wire \heichips25_sap3/_0521_ ;
 wire \heichips25_sap3/_0522_ ;
 wire \heichips25_sap3/_0523_ ;
 wire \heichips25_sap3/_0524_ ;
 wire \heichips25_sap3/_0525_ ;
 wire \heichips25_sap3/_0526_ ;
 wire \heichips25_sap3/_0527_ ;
 wire \heichips25_sap3/_0528_ ;
 wire \heichips25_sap3/_0529_ ;
 wire \heichips25_sap3/_0530_ ;
 wire \heichips25_sap3/_0531_ ;
 wire \heichips25_sap3/_0532_ ;
 wire \heichips25_sap3/_0533_ ;
 wire \heichips25_sap3/_0534_ ;
 wire \heichips25_sap3/_0535_ ;
 wire \heichips25_sap3/_0536_ ;
 wire \heichips25_sap3/_0537_ ;
 wire \heichips25_sap3/_0538_ ;
 wire \heichips25_sap3/_0539_ ;
 wire \heichips25_sap3/_0540_ ;
 wire \heichips25_sap3/_0541_ ;
 wire \heichips25_sap3/_0542_ ;
 wire \heichips25_sap3/_0543_ ;
 wire \heichips25_sap3/_0544_ ;
 wire \heichips25_sap3/_0545_ ;
 wire \heichips25_sap3/_0546_ ;
 wire \heichips25_sap3/_0547_ ;
 wire \heichips25_sap3/_0548_ ;
 wire \heichips25_sap3/_0549_ ;
 wire \heichips25_sap3/_0550_ ;
 wire \heichips25_sap3/_0551_ ;
 wire \heichips25_sap3/_0552_ ;
 wire \heichips25_sap3/_0553_ ;
 wire \heichips25_sap3/_0554_ ;
 wire \heichips25_sap3/_0555_ ;
 wire \heichips25_sap3/_0556_ ;
 wire \heichips25_sap3/_0557_ ;
 wire \heichips25_sap3/_0558_ ;
 wire \heichips25_sap3/_0559_ ;
 wire \heichips25_sap3/_0560_ ;
 wire \heichips25_sap3/_0561_ ;
 wire \heichips25_sap3/_0562_ ;
 wire \heichips25_sap3/_0563_ ;
 wire \heichips25_sap3/_0564_ ;
 wire \heichips25_sap3/_0565_ ;
 wire \heichips25_sap3/_0566_ ;
 wire \heichips25_sap3/_0567_ ;
 wire \heichips25_sap3/_0568_ ;
 wire \heichips25_sap3/_0569_ ;
 wire \heichips25_sap3/_0570_ ;
 wire \heichips25_sap3/_0571_ ;
 wire \heichips25_sap3/_0572_ ;
 wire \heichips25_sap3/_0573_ ;
 wire \heichips25_sap3/_0574_ ;
 wire \heichips25_sap3/_0575_ ;
 wire \heichips25_sap3/_0576_ ;
 wire \heichips25_sap3/_0577_ ;
 wire \heichips25_sap3/_0578_ ;
 wire \heichips25_sap3/_0579_ ;
 wire \heichips25_sap3/_0580_ ;
 wire \heichips25_sap3/_0581_ ;
 wire \heichips25_sap3/_0582_ ;
 wire \heichips25_sap3/_0583_ ;
 wire \heichips25_sap3/_0584_ ;
 wire \heichips25_sap3/_0585_ ;
 wire \heichips25_sap3/_0586_ ;
 wire \heichips25_sap3/_0587_ ;
 wire \heichips25_sap3/_0588_ ;
 wire \heichips25_sap3/_0589_ ;
 wire \heichips25_sap3/_0590_ ;
 wire \heichips25_sap3/_0591_ ;
 wire \heichips25_sap3/_0592_ ;
 wire \heichips25_sap3/_0593_ ;
 wire \heichips25_sap3/_0594_ ;
 wire \heichips25_sap3/_0595_ ;
 wire \heichips25_sap3/_0596_ ;
 wire \heichips25_sap3/_0597_ ;
 wire \heichips25_sap3/_0598_ ;
 wire \heichips25_sap3/_0599_ ;
 wire \heichips25_sap3/_0600_ ;
 wire \heichips25_sap3/_0601_ ;
 wire \heichips25_sap3/_0602_ ;
 wire \heichips25_sap3/_0603_ ;
 wire \heichips25_sap3/_0604_ ;
 wire \heichips25_sap3/_0605_ ;
 wire \heichips25_sap3/_0606_ ;
 wire \heichips25_sap3/_0607_ ;
 wire \heichips25_sap3/_0608_ ;
 wire \heichips25_sap3/_0609_ ;
 wire \heichips25_sap3/_0610_ ;
 wire \heichips25_sap3/_0611_ ;
 wire \heichips25_sap3/_0612_ ;
 wire \heichips25_sap3/_0613_ ;
 wire \heichips25_sap3/_0614_ ;
 wire \heichips25_sap3/_0615_ ;
 wire \heichips25_sap3/_0616_ ;
 wire \heichips25_sap3/_0617_ ;
 wire \heichips25_sap3/_0618_ ;
 wire \heichips25_sap3/_0619_ ;
 wire \heichips25_sap3/_0620_ ;
 wire \heichips25_sap3/_0621_ ;
 wire \heichips25_sap3/_0622_ ;
 wire \heichips25_sap3/_0623_ ;
 wire \heichips25_sap3/_0624_ ;
 wire \heichips25_sap3/_0625_ ;
 wire \heichips25_sap3/_0626_ ;
 wire \heichips25_sap3/_0627_ ;
 wire \heichips25_sap3/_0628_ ;
 wire \heichips25_sap3/_0629_ ;
 wire \heichips25_sap3/_0630_ ;
 wire \heichips25_sap3/_0631_ ;
 wire \heichips25_sap3/_0632_ ;
 wire \heichips25_sap3/_0633_ ;
 wire \heichips25_sap3/_0634_ ;
 wire \heichips25_sap3/_0635_ ;
 wire \heichips25_sap3/_0636_ ;
 wire \heichips25_sap3/_0637_ ;
 wire \heichips25_sap3/_0638_ ;
 wire \heichips25_sap3/_0639_ ;
 wire \heichips25_sap3/_0640_ ;
 wire \heichips25_sap3/_0641_ ;
 wire \heichips25_sap3/_0642_ ;
 wire \heichips25_sap3/_0643_ ;
 wire \heichips25_sap3/_0644_ ;
 wire \heichips25_sap3/_0645_ ;
 wire \heichips25_sap3/_0646_ ;
 wire \heichips25_sap3/_0647_ ;
 wire \heichips25_sap3/_0648_ ;
 wire \heichips25_sap3/_0649_ ;
 wire \heichips25_sap3/_0650_ ;
 wire \heichips25_sap3/_0651_ ;
 wire \heichips25_sap3/_0652_ ;
 wire \heichips25_sap3/_0653_ ;
 wire \heichips25_sap3/_0654_ ;
 wire \heichips25_sap3/_0655_ ;
 wire \heichips25_sap3/_0656_ ;
 wire \heichips25_sap3/_0657_ ;
 wire \heichips25_sap3/_0658_ ;
 wire \heichips25_sap3/_0659_ ;
 wire \heichips25_sap3/_0660_ ;
 wire \heichips25_sap3/_0661_ ;
 wire \heichips25_sap3/_0662_ ;
 wire \heichips25_sap3/_0663_ ;
 wire \heichips25_sap3/_0664_ ;
 wire \heichips25_sap3/_0665_ ;
 wire \heichips25_sap3/_0666_ ;
 wire \heichips25_sap3/_0667_ ;
 wire \heichips25_sap3/_0668_ ;
 wire \heichips25_sap3/_0669_ ;
 wire \heichips25_sap3/_0670_ ;
 wire \heichips25_sap3/_0671_ ;
 wire \heichips25_sap3/_0672_ ;
 wire \heichips25_sap3/_0673_ ;
 wire \heichips25_sap3/_0674_ ;
 wire \heichips25_sap3/_0675_ ;
 wire \heichips25_sap3/_0676_ ;
 wire \heichips25_sap3/_0677_ ;
 wire \heichips25_sap3/_0678_ ;
 wire \heichips25_sap3/_0679_ ;
 wire \heichips25_sap3/_0680_ ;
 wire \heichips25_sap3/_0681_ ;
 wire \heichips25_sap3/_0682_ ;
 wire \heichips25_sap3/_0683_ ;
 wire \heichips25_sap3/_0684_ ;
 wire \heichips25_sap3/_0685_ ;
 wire \heichips25_sap3/_0686_ ;
 wire \heichips25_sap3/_0687_ ;
 wire \heichips25_sap3/_0688_ ;
 wire \heichips25_sap3/_0689_ ;
 wire \heichips25_sap3/_0690_ ;
 wire \heichips25_sap3/_0691_ ;
 wire \heichips25_sap3/_0692_ ;
 wire \heichips25_sap3/_0693_ ;
 wire \heichips25_sap3/_0694_ ;
 wire \heichips25_sap3/_0695_ ;
 wire \heichips25_sap3/_0696_ ;
 wire \heichips25_sap3/_0697_ ;
 wire \heichips25_sap3/_0698_ ;
 wire \heichips25_sap3/_0699_ ;
 wire \heichips25_sap3/_0700_ ;
 wire \heichips25_sap3/_0701_ ;
 wire \heichips25_sap3/_0702_ ;
 wire \heichips25_sap3/_0703_ ;
 wire \heichips25_sap3/_0704_ ;
 wire \heichips25_sap3/_0705_ ;
 wire \heichips25_sap3/_0706_ ;
 wire \heichips25_sap3/_0707_ ;
 wire \heichips25_sap3/_0708_ ;
 wire \heichips25_sap3/_0709_ ;
 wire \heichips25_sap3/_0710_ ;
 wire \heichips25_sap3/_0711_ ;
 wire \heichips25_sap3/_0712_ ;
 wire \heichips25_sap3/_0713_ ;
 wire \heichips25_sap3/_0714_ ;
 wire \heichips25_sap3/_0715_ ;
 wire \heichips25_sap3/_0716_ ;
 wire \heichips25_sap3/_0717_ ;
 wire \heichips25_sap3/_0718_ ;
 wire \heichips25_sap3/_0719_ ;
 wire \heichips25_sap3/_0720_ ;
 wire \heichips25_sap3/_0721_ ;
 wire \heichips25_sap3/_0722_ ;
 wire \heichips25_sap3/_0723_ ;
 wire \heichips25_sap3/_0724_ ;
 wire \heichips25_sap3/_0725_ ;
 wire \heichips25_sap3/_0726_ ;
 wire \heichips25_sap3/_0727_ ;
 wire \heichips25_sap3/_0728_ ;
 wire \heichips25_sap3/_0729_ ;
 wire \heichips25_sap3/_0730_ ;
 wire \heichips25_sap3/_0731_ ;
 wire \heichips25_sap3/_0732_ ;
 wire \heichips25_sap3/_0733_ ;
 wire \heichips25_sap3/_0734_ ;
 wire \heichips25_sap3/_0735_ ;
 wire \heichips25_sap3/_0736_ ;
 wire \heichips25_sap3/_0737_ ;
 wire \heichips25_sap3/_0738_ ;
 wire \heichips25_sap3/_0739_ ;
 wire \heichips25_sap3/_0740_ ;
 wire \heichips25_sap3/_0741_ ;
 wire \heichips25_sap3/_0742_ ;
 wire \heichips25_sap3/_0743_ ;
 wire \heichips25_sap3/_0744_ ;
 wire \heichips25_sap3/_0745_ ;
 wire \heichips25_sap3/_0746_ ;
 wire \heichips25_sap3/_0747_ ;
 wire \heichips25_sap3/_0748_ ;
 wire \heichips25_sap3/_0749_ ;
 wire \heichips25_sap3/_0750_ ;
 wire \heichips25_sap3/_0751_ ;
 wire \heichips25_sap3/_0752_ ;
 wire \heichips25_sap3/_0753_ ;
 wire \heichips25_sap3/_0754_ ;
 wire \heichips25_sap3/_0755_ ;
 wire \heichips25_sap3/_0756_ ;
 wire \heichips25_sap3/_0757_ ;
 wire \heichips25_sap3/_0758_ ;
 wire \heichips25_sap3/_0759_ ;
 wire \heichips25_sap3/_0760_ ;
 wire \heichips25_sap3/_0761_ ;
 wire \heichips25_sap3/_0762_ ;
 wire \heichips25_sap3/_0763_ ;
 wire \heichips25_sap3/_0764_ ;
 wire \heichips25_sap3/_0765_ ;
 wire \heichips25_sap3/_0766_ ;
 wire \heichips25_sap3/_0767_ ;
 wire \heichips25_sap3/_0768_ ;
 wire \heichips25_sap3/_0769_ ;
 wire \heichips25_sap3/_0770_ ;
 wire \heichips25_sap3/_0771_ ;
 wire \heichips25_sap3/_0772_ ;
 wire \heichips25_sap3/_0773_ ;
 wire \heichips25_sap3/_0774_ ;
 wire \heichips25_sap3/_0775_ ;
 wire \heichips25_sap3/_0776_ ;
 wire \heichips25_sap3/_0777_ ;
 wire \heichips25_sap3/_0778_ ;
 wire \heichips25_sap3/_0779_ ;
 wire \heichips25_sap3/_0780_ ;
 wire \heichips25_sap3/_0781_ ;
 wire \heichips25_sap3/_0782_ ;
 wire \heichips25_sap3/_0783_ ;
 wire \heichips25_sap3/_0784_ ;
 wire \heichips25_sap3/_0785_ ;
 wire \heichips25_sap3/_0786_ ;
 wire \heichips25_sap3/_0787_ ;
 wire \heichips25_sap3/_0788_ ;
 wire \heichips25_sap3/_0789_ ;
 wire \heichips25_sap3/_0790_ ;
 wire \heichips25_sap3/_0791_ ;
 wire \heichips25_sap3/_0792_ ;
 wire \heichips25_sap3/_0793_ ;
 wire \heichips25_sap3/_0794_ ;
 wire \heichips25_sap3/_0795_ ;
 wire \heichips25_sap3/_0796_ ;
 wire \heichips25_sap3/_0797_ ;
 wire \heichips25_sap3/_0798_ ;
 wire \heichips25_sap3/_0799_ ;
 wire \heichips25_sap3/_0800_ ;
 wire \heichips25_sap3/_0801_ ;
 wire \heichips25_sap3/_0802_ ;
 wire \heichips25_sap3/_0803_ ;
 wire \heichips25_sap3/_0804_ ;
 wire \heichips25_sap3/_0805_ ;
 wire \heichips25_sap3/_0806_ ;
 wire \heichips25_sap3/_0807_ ;
 wire \heichips25_sap3/_0808_ ;
 wire \heichips25_sap3/_0809_ ;
 wire \heichips25_sap3/_0810_ ;
 wire \heichips25_sap3/_0811_ ;
 wire \heichips25_sap3/_0812_ ;
 wire \heichips25_sap3/_0813_ ;
 wire \heichips25_sap3/_0814_ ;
 wire \heichips25_sap3/_0815_ ;
 wire \heichips25_sap3/_0816_ ;
 wire \heichips25_sap3/_0817_ ;
 wire \heichips25_sap3/_0818_ ;
 wire \heichips25_sap3/_0819_ ;
 wire \heichips25_sap3/_0820_ ;
 wire \heichips25_sap3/_0821_ ;
 wire \heichips25_sap3/_0822_ ;
 wire \heichips25_sap3/_0823_ ;
 wire \heichips25_sap3/_0824_ ;
 wire \heichips25_sap3/_0825_ ;
 wire \heichips25_sap3/_0826_ ;
 wire \heichips25_sap3/_0827_ ;
 wire \heichips25_sap3/_0828_ ;
 wire \heichips25_sap3/_0829_ ;
 wire \heichips25_sap3/_0830_ ;
 wire \heichips25_sap3/_0831_ ;
 wire \heichips25_sap3/_0832_ ;
 wire \heichips25_sap3/_0833_ ;
 wire \heichips25_sap3/_0834_ ;
 wire \heichips25_sap3/_0835_ ;
 wire \heichips25_sap3/_0836_ ;
 wire \heichips25_sap3/_0837_ ;
 wire \heichips25_sap3/_0838_ ;
 wire \heichips25_sap3/_0839_ ;
 wire \heichips25_sap3/_0840_ ;
 wire \heichips25_sap3/_0841_ ;
 wire \heichips25_sap3/_0842_ ;
 wire \heichips25_sap3/_0843_ ;
 wire \heichips25_sap3/_0844_ ;
 wire \heichips25_sap3/_0845_ ;
 wire \heichips25_sap3/_0846_ ;
 wire \heichips25_sap3/_0847_ ;
 wire \heichips25_sap3/_0848_ ;
 wire \heichips25_sap3/_0849_ ;
 wire \heichips25_sap3/_0850_ ;
 wire \heichips25_sap3/_0851_ ;
 wire \heichips25_sap3/_0852_ ;
 wire \heichips25_sap3/_0853_ ;
 wire \heichips25_sap3/_0854_ ;
 wire \heichips25_sap3/_0855_ ;
 wire \heichips25_sap3/_0856_ ;
 wire \heichips25_sap3/_0857_ ;
 wire \heichips25_sap3/_0858_ ;
 wire \heichips25_sap3/_0859_ ;
 wire \heichips25_sap3/_0860_ ;
 wire \heichips25_sap3/_0861_ ;
 wire \heichips25_sap3/_0862_ ;
 wire \heichips25_sap3/_0863_ ;
 wire \heichips25_sap3/_0864_ ;
 wire \heichips25_sap3/_0865_ ;
 wire \heichips25_sap3/_0866_ ;
 wire \heichips25_sap3/_0867_ ;
 wire \heichips25_sap3/_0868_ ;
 wire \heichips25_sap3/_0869_ ;
 wire \heichips25_sap3/_0870_ ;
 wire \heichips25_sap3/_0871_ ;
 wire \heichips25_sap3/_0872_ ;
 wire \heichips25_sap3/_0873_ ;
 wire \heichips25_sap3/_0874_ ;
 wire \heichips25_sap3/_0875_ ;
 wire \heichips25_sap3/_0876_ ;
 wire \heichips25_sap3/_0877_ ;
 wire \heichips25_sap3/_0878_ ;
 wire \heichips25_sap3/_0879_ ;
 wire \heichips25_sap3/_0880_ ;
 wire \heichips25_sap3/_0881_ ;
 wire \heichips25_sap3/_0882_ ;
 wire \heichips25_sap3/_0883_ ;
 wire \heichips25_sap3/_0884_ ;
 wire \heichips25_sap3/_0885_ ;
 wire \heichips25_sap3/_0886_ ;
 wire \heichips25_sap3/_0887_ ;
 wire \heichips25_sap3/_0888_ ;
 wire \heichips25_sap3/_0889_ ;
 wire \heichips25_sap3/_0890_ ;
 wire \heichips25_sap3/_0891_ ;
 wire \heichips25_sap3/_0892_ ;
 wire \heichips25_sap3/_0893_ ;
 wire \heichips25_sap3/_0894_ ;
 wire \heichips25_sap3/_0895_ ;
 wire \heichips25_sap3/_0896_ ;
 wire \heichips25_sap3/_0897_ ;
 wire \heichips25_sap3/_0898_ ;
 wire \heichips25_sap3/_0899_ ;
 wire \heichips25_sap3/_0900_ ;
 wire \heichips25_sap3/_0901_ ;
 wire \heichips25_sap3/_0902_ ;
 wire \heichips25_sap3/_0903_ ;
 wire \heichips25_sap3/_0904_ ;
 wire \heichips25_sap3/_0905_ ;
 wire \heichips25_sap3/_0906_ ;
 wire \heichips25_sap3/_0907_ ;
 wire \heichips25_sap3/_0908_ ;
 wire \heichips25_sap3/_0909_ ;
 wire \heichips25_sap3/_0910_ ;
 wire \heichips25_sap3/_0911_ ;
 wire \heichips25_sap3/_0912_ ;
 wire \heichips25_sap3/_0913_ ;
 wire \heichips25_sap3/_0914_ ;
 wire \heichips25_sap3/_0915_ ;
 wire \heichips25_sap3/_0916_ ;
 wire \heichips25_sap3/_0917_ ;
 wire \heichips25_sap3/_0918_ ;
 wire \heichips25_sap3/_0919_ ;
 wire \heichips25_sap3/_0920_ ;
 wire \heichips25_sap3/_0921_ ;
 wire \heichips25_sap3/_0922_ ;
 wire \heichips25_sap3/_0923_ ;
 wire \heichips25_sap3/_0924_ ;
 wire \heichips25_sap3/_0925_ ;
 wire \heichips25_sap3/_0926_ ;
 wire \heichips25_sap3/_0927_ ;
 wire \heichips25_sap3/_0928_ ;
 wire \heichips25_sap3/_0929_ ;
 wire \heichips25_sap3/_0930_ ;
 wire \heichips25_sap3/_0931_ ;
 wire \heichips25_sap3/_0932_ ;
 wire \heichips25_sap3/_0933_ ;
 wire \heichips25_sap3/_0934_ ;
 wire \heichips25_sap3/_0935_ ;
 wire \heichips25_sap3/_0936_ ;
 wire \heichips25_sap3/_0937_ ;
 wire \heichips25_sap3/_0938_ ;
 wire \heichips25_sap3/_0939_ ;
 wire \heichips25_sap3/_0940_ ;
 wire \heichips25_sap3/_0941_ ;
 wire \heichips25_sap3/_0942_ ;
 wire \heichips25_sap3/_0943_ ;
 wire \heichips25_sap3/_0944_ ;
 wire \heichips25_sap3/_0945_ ;
 wire \heichips25_sap3/_0946_ ;
 wire \heichips25_sap3/_0947_ ;
 wire \heichips25_sap3/_0948_ ;
 wire \heichips25_sap3/_0949_ ;
 wire \heichips25_sap3/_0950_ ;
 wire \heichips25_sap3/_0951_ ;
 wire \heichips25_sap3/_0952_ ;
 wire \heichips25_sap3/_0953_ ;
 wire \heichips25_sap3/_0954_ ;
 wire \heichips25_sap3/_0955_ ;
 wire \heichips25_sap3/_0956_ ;
 wire \heichips25_sap3/_0957_ ;
 wire \heichips25_sap3/_0958_ ;
 wire \heichips25_sap3/_0959_ ;
 wire \heichips25_sap3/_0960_ ;
 wire \heichips25_sap3/_0961_ ;
 wire \heichips25_sap3/_0962_ ;
 wire \heichips25_sap3/_0963_ ;
 wire \heichips25_sap3/_0964_ ;
 wire \heichips25_sap3/_0965_ ;
 wire \heichips25_sap3/_0966_ ;
 wire \heichips25_sap3/_0967_ ;
 wire \heichips25_sap3/_0968_ ;
 wire \heichips25_sap3/_0969_ ;
 wire \heichips25_sap3/_0970_ ;
 wire \heichips25_sap3/_0971_ ;
 wire \heichips25_sap3/_0972_ ;
 wire \heichips25_sap3/_0973_ ;
 wire \heichips25_sap3/_0974_ ;
 wire \heichips25_sap3/_0975_ ;
 wire \heichips25_sap3/_0976_ ;
 wire \heichips25_sap3/_0977_ ;
 wire \heichips25_sap3/_0978_ ;
 wire \heichips25_sap3/_0979_ ;
 wire \heichips25_sap3/_0980_ ;
 wire \heichips25_sap3/_0981_ ;
 wire \heichips25_sap3/_0982_ ;
 wire \heichips25_sap3/_0983_ ;
 wire \heichips25_sap3/_0984_ ;
 wire \heichips25_sap3/_0985_ ;
 wire \heichips25_sap3/_0986_ ;
 wire \heichips25_sap3/_0987_ ;
 wire \heichips25_sap3/_0988_ ;
 wire \heichips25_sap3/_0989_ ;
 wire \heichips25_sap3/_0990_ ;
 wire \heichips25_sap3/_0991_ ;
 wire \heichips25_sap3/_0992_ ;
 wire \heichips25_sap3/_0993_ ;
 wire \heichips25_sap3/_0994_ ;
 wire \heichips25_sap3/_0995_ ;
 wire \heichips25_sap3/_0996_ ;
 wire \heichips25_sap3/_0997_ ;
 wire \heichips25_sap3/_0998_ ;
 wire \heichips25_sap3/_0999_ ;
 wire \heichips25_sap3/_1000_ ;
 wire \heichips25_sap3/_1001_ ;
 wire \heichips25_sap3/_1002_ ;
 wire \heichips25_sap3/_1003_ ;
 wire \heichips25_sap3/_1004_ ;
 wire \heichips25_sap3/_1005_ ;
 wire \heichips25_sap3/_1006_ ;
 wire \heichips25_sap3/_1007_ ;
 wire \heichips25_sap3/_1008_ ;
 wire \heichips25_sap3/_1009_ ;
 wire \heichips25_sap3/_1010_ ;
 wire \heichips25_sap3/_1011_ ;
 wire \heichips25_sap3/_1012_ ;
 wire \heichips25_sap3/_1013_ ;
 wire \heichips25_sap3/_1014_ ;
 wire \heichips25_sap3/_1015_ ;
 wire \heichips25_sap3/_1016_ ;
 wire \heichips25_sap3/_1017_ ;
 wire \heichips25_sap3/_1018_ ;
 wire \heichips25_sap3/_1019_ ;
 wire \heichips25_sap3/_1020_ ;
 wire \heichips25_sap3/_1021_ ;
 wire \heichips25_sap3/_1022_ ;
 wire \heichips25_sap3/_1023_ ;
 wire \heichips25_sap3/_1024_ ;
 wire \heichips25_sap3/_1025_ ;
 wire \heichips25_sap3/_1026_ ;
 wire \heichips25_sap3/_1027_ ;
 wire \heichips25_sap3/_1028_ ;
 wire \heichips25_sap3/_1029_ ;
 wire \heichips25_sap3/_1030_ ;
 wire \heichips25_sap3/_1031_ ;
 wire \heichips25_sap3/_1032_ ;
 wire \heichips25_sap3/_1033_ ;
 wire \heichips25_sap3/_1034_ ;
 wire \heichips25_sap3/_1035_ ;
 wire \heichips25_sap3/_1036_ ;
 wire \heichips25_sap3/_1037_ ;
 wire \heichips25_sap3/_1038_ ;
 wire \heichips25_sap3/_1039_ ;
 wire \heichips25_sap3/_1040_ ;
 wire \heichips25_sap3/_1041_ ;
 wire \heichips25_sap3/_1042_ ;
 wire \heichips25_sap3/_1043_ ;
 wire \heichips25_sap3/_1044_ ;
 wire \heichips25_sap3/_1045_ ;
 wire \heichips25_sap3/_1046_ ;
 wire \heichips25_sap3/_1047_ ;
 wire \heichips25_sap3/_1048_ ;
 wire \heichips25_sap3/_1049_ ;
 wire \heichips25_sap3/_1050_ ;
 wire \heichips25_sap3/_1051_ ;
 wire \heichips25_sap3/_1052_ ;
 wire \heichips25_sap3/_1053_ ;
 wire \heichips25_sap3/_1054_ ;
 wire \heichips25_sap3/_1055_ ;
 wire \heichips25_sap3/_1056_ ;
 wire \heichips25_sap3/_1057_ ;
 wire \heichips25_sap3/_1058_ ;
 wire \heichips25_sap3/_1059_ ;
 wire \heichips25_sap3/_1060_ ;
 wire \heichips25_sap3/_1061_ ;
 wire \heichips25_sap3/_1062_ ;
 wire \heichips25_sap3/_1063_ ;
 wire \heichips25_sap3/_1064_ ;
 wire \heichips25_sap3/_1065_ ;
 wire \heichips25_sap3/_1066_ ;
 wire \heichips25_sap3/_1067_ ;
 wire \heichips25_sap3/_1068_ ;
 wire \heichips25_sap3/_1069_ ;
 wire \heichips25_sap3/_1070_ ;
 wire \heichips25_sap3/_1071_ ;
 wire \heichips25_sap3/_1072_ ;
 wire \heichips25_sap3/_1073_ ;
 wire \heichips25_sap3/_1074_ ;
 wire \heichips25_sap3/_1075_ ;
 wire \heichips25_sap3/_1076_ ;
 wire \heichips25_sap3/_1077_ ;
 wire \heichips25_sap3/_1078_ ;
 wire \heichips25_sap3/_1079_ ;
 wire \heichips25_sap3/_1080_ ;
 wire \heichips25_sap3/_1081_ ;
 wire \heichips25_sap3/_1082_ ;
 wire \heichips25_sap3/_1083_ ;
 wire \heichips25_sap3/_1084_ ;
 wire \heichips25_sap3/_1085_ ;
 wire \heichips25_sap3/_1086_ ;
 wire \heichips25_sap3/_1087_ ;
 wire \heichips25_sap3/_1088_ ;
 wire \heichips25_sap3/_1089_ ;
 wire \heichips25_sap3/_1090_ ;
 wire \heichips25_sap3/_1091_ ;
 wire \heichips25_sap3/_1092_ ;
 wire \heichips25_sap3/_1093_ ;
 wire \heichips25_sap3/_1094_ ;
 wire \heichips25_sap3/_1095_ ;
 wire \heichips25_sap3/_1096_ ;
 wire \heichips25_sap3/_1097_ ;
 wire \heichips25_sap3/_1098_ ;
 wire \heichips25_sap3/_1099_ ;
 wire \heichips25_sap3/_1100_ ;
 wire \heichips25_sap3/_1101_ ;
 wire \heichips25_sap3/_1102_ ;
 wire \heichips25_sap3/_1103_ ;
 wire \heichips25_sap3/_1104_ ;
 wire \heichips25_sap3/_1105_ ;
 wire \heichips25_sap3/_1106_ ;
 wire \heichips25_sap3/_1107_ ;
 wire \heichips25_sap3/_1108_ ;
 wire \heichips25_sap3/_1109_ ;
 wire \heichips25_sap3/_1110_ ;
 wire \heichips25_sap3/_1111_ ;
 wire \heichips25_sap3/_1112_ ;
 wire \heichips25_sap3/_1113_ ;
 wire \heichips25_sap3/_1114_ ;
 wire \heichips25_sap3/_1115_ ;
 wire \heichips25_sap3/_1116_ ;
 wire \heichips25_sap3/_1117_ ;
 wire \heichips25_sap3/_1118_ ;
 wire \heichips25_sap3/_1119_ ;
 wire \heichips25_sap3/_1120_ ;
 wire \heichips25_sap3/_1121_ ;
 wire \heichips25_sap3/_1122_ ;
 wire \heichips25_sap3/_1123_ ;
 wire \heichips25_sap3/_1124_ ;
 wire \heichips25_sap3/_1125_ ;
 wire \heichips25_sap3/_1126_ ;
 wire \heichips25_sap3/_1127_ ;
 wire \heichips25_sap3/_1128_ ;
 wire \heichips25_sap3/_1129_ ;
 wire \heichips25_sap3/_1130_ ;
 wire \heichips25_sap3/_1131_ ;
 wire \heichips25_sap3/_1132_ ;
 wire \heichips25_sap3/_1133_ ;
 wire \heichips25_sap3/_1134_ ;
 wire \heichips25_sap3/_1135_ ;
 wire \heichips25_sap3/_1136_ ;
 wire \heichips25_sap3/_1137_ ;
 wire \heichips25_sap3/_1138_ ;
 wire \heichips25_sap3/_1139_ ;
 wire \heichips25_sap3/_1140_ ;
 wire \heichips25_sap3/_1141_ ;
 wire \heichips25_sap3/_1142_ ;
 wire \heichips25_sap3/_1143_ ;
 wire \heichips25_sap3/_1144_ ;
 wire \heichips25_sap3/_1145_ ;
 wire \heichips25_sap3/_1146_ ;
 wire \heichips25_sap3/_1147_ ;
 wire \heichips25_sap3/_1148_ ;
 wire \heichips25_sap3/_1149_ ;
 wire \heichips25_sap3/_1150_ ;
 wire \heichips25_sap3/_1151_ ;
 wire \heichips25_sap3/_1152_ ;
 wire \heichips25_sap3/_1153_ ;
 wire \heichips25_sap3/_1154_ ;
 wire \heichips25_sap3/_1155_ ;
 wire \heichips25_sap3/_1156_ ;
 wire \heichips25_sap3/_1157_ ;
 wire \heichips25_sap3/_1158_ ;
 wire \heichips25_sap3/_1159_ ;
 wire \heichips25_sap3/_1160_ ;
 wire \heichips25_sap3/_1161_ ;
 wire \heichips25_sap3/_1162_ ;
 wire \heichips25_sap3/_1163_ ;
 wire \heichips25_sap3/_1164_ ;
 wire \heichips25_sap3/_1165_ ;
 wire \heichips25_sap3/_1166_ ;
 wire \heichips25_sap3/_1167_ ;
 wire \heichips25_sap3/_1168_ ;
 wire \heichips25_sap3/_1169_ ;
 wire \heichips25_sap3/_1170_ ;
 wire \heichips25_sap3/_1171_ ;
 wire \heichips25_sap3/_1172_ ;
 wire \heichips25_sap3/_1173_ ;
 wire \heichips25_sap3/_1174_ ;
 wire \heichips25_sap3/_1175_ ;
 wire \heichips25_sap3/_1176_ ;
 wire \heichips25_sap3/_1177_ ;
 wire \heichips25_sap3/_1178_ ;
 wire \heichips25_sap3/_1179_ ;
 wire \heichips25_sap3/_1180_ ;
 wire \heichips25_sap3/_1181_ ;
 wire \heichips25_sap3/_1182_ ;
 wire \heichips25_sap3/_1183_ ;
 wire \heichips25_sap3/_1184_ ;
 wire \heichips25_sap3/_1185_ ;
 wire \heichips25_sap3/_1186_ ;
 wire \heichips25_sap3/_1187_ ;
 wire \heichips25_sap3/_1188_ ;
 wire \heichips25_sap3/_1189_ ;
 wire \heichips25_sap3/_1190_ ;
 wire \heichips25_sap3/_1191_ ;
 wire \heichips25_sap3/_1192_ ;
 wire \heichips25_sap3/_1193_ ;
 wire \heichips25_sap3/_1194_ ;
 wire \heichips25_sap3/_1195_ ;
 wire \heichips25_sap3/_1196_ ;
 wire \heichips25_sap3/_1197_ ;
 wire \heichips25_sap3/_1198_ ;
 wire \heichips25_sap3/_1199_ ;
 wire \heichips25_sap3/_1200_ ;
 wire \heichips25_sap3/_1201_ ;
 wire \heichips25_sap3/_1202_ ;
 wire \heichips25_sap3/_1203_ ;
 wire \heichips25_sap3/_1204_ ;
 wire \heichips25_sap3/_1205_ ;
 wire \heichips25_sap3/_1206_ ;
 wire \heichips25_sap3/_1207_ ;
 wire \heichips25_sap3/_1208_ ;
 wire \heichips25_sap3/_1209_ ;
 wire \heichips25_sap3/_1210_ ;
 wire \heichips25_sap3/_1211_ ;
 wire \heichips25_sap3/_1212_ ;
 wire \heichips25_sap3/_1213_ ;
 wire \heichips25_sap3/_1214_ ;
 wire \heichips25_sap3/_1215_ ;
 wire \heichips25_sap3/_1216_ ;
 wire \heichips25_sap3/_1217_ ;
 wire \heichips25_sap3/_1218_ ;
 wire \heichips25_sap3/_1219_ ;
 wire \heichips25_sap3/_1220_ ;
 wire \heichips25_sap3/_1221_ ;
 wire \heichips25_sap3/_1222_ ;
 wire \heichips25_sap3/_1223_ ;
 wire \heichips25_sap3/_1224_ ;
 wire \heichips25_sap3/_1225_ ;
 wire \heichips25_sap3/_1226_ ;
 wire \heichips25_sap3/_1227_ ;
 wire \heichips25_sap3/_1228_ ;
 wire \heichips25_sap3/_1229_ ;
 wire \heichips25_sap3/_1230_ ;
 wire \heichips25_sap3/_1231_ ;
 wire \heichips25_sap3/_1232_ ;
 wire \heichips25_sap3/_1233_ ;
 wire \heichips25_sap3/_1234_ ;
 wire \heichips25_sap3/_1235_ ;
 wire \heichips25_sap3/_1236_ ;
 wire \heichips25_sap3/_1237_ ;
 wire \heichips25_sap3/_1238_ ;
 wire \heichips25_sap3/_1239_ ;
 wire \heichips25_sap3/_1240_ ;
 wire \heichips25_sap3/_1241_ ;
 wire \heichips25_sap3/_1242_ ;
 wire \heichips25_sap3/_1243_ ;
 wire \heichips25_sap3/_1244_ ;
 wire \heichips25_sap3/_1245_ ;
 wire \heichips25_sap3/_1246_ ;
 wire \heichips25_sap3/_1247_ ;
 wire \heichips25_sap3/_1248_ ;
 wire \heichips25_sap3/_1249_ ;
 wire \heichips25_sap3/_1250_ ;
 wire \heichips25_sap3/_1251_ ;
 wire \heichips25_sap3/_1252_ ;
 wire \heichips25_sap3/_1253_ ;
 wire \heichips25_sap3/_1254_ ;
 wire \heichips25_sap3/_1255_ ;
 wire \heichips25_sap3/_1256_ ;
 wire \heichips25_sap3/_1257_ ;
 wire \heichips25_sap3/_1258_ ;
 wire \heichips25_sap3/_1259_ ;
 wire \heichips25_sap3/_1260_ ;
 wire \heichips25_sap3/_1261_ ;
 wire \heichips25_sap3/_1262_ ;
 wire \heichips25_sap3/_1263_ ;
 wire \heichips25_sap3/_1264_ ;
 wire \heichips25_sap3/_1265_ ;
 wire \heichips25_sap3/_1266_ ;
 wire \heichips25_sap3/_1267_ ;
 wire \heichips25_sap3/_1268_ ;
 wire \heichips25_sap3/_1269_ ;
 wire \heichips25_sap3/_1270_ ;
 wire \heichips25_sap3/_1271_ ;
 wire \heichips25_sap3/_1272_ ;
 wire \heichips25_sap3/_1273_ ;
 wire \heichips25_sap3/_1274_ ;
 wire \heichips25_sap3/_1275_ ;
 wire \heichips25_sap3/_1276_ ;
 wire \heichips25_sap3/_1277_ ;
 wire \heichips25_sap3/_1278_ ;
 wire \heichips25_sap3/_1279_ ;
 wire \heichips25_sap3/_1280_ ;
 wire \heichips25_sap3/_1281_ ;
 wire \heichips25_sap3/_1282_ ;
 wire \heichips25_sap3/_1283_ ;
 wire \heichips25_sap3/_1284_ ;
 wire \heichips25_sap3/_1285_ ;
 wire \heichips25_sap3/_1286_ ;
 wire \heichips25_sap3/_1287_ ;
 wire \heichips25_sap3/_1288_ ;
 wire \heichips25_sap3/_1289_ ;
 wire \heichips25_sap3/_1290_ ;
 wire \heichips25_sap3/_1291_ ;
 wire \heichips25_sap3/_1292_ ;
 wire \heichips25_sap3/_1293_ ;
 wire \heichips25_sap3/_1294_ ;
 wire \heichips25_sap3/_1295_ ;
 wire \heichips25_sap3/_1296_ ;
 wire \heichips25_sap3/_1297_ ;
 wire \heichips25_sap3/_1298_ ;
 wire \heichips25_sap3/_1299_ ;
 wire \heichips25_sap3/_1300_ ;
 wire \heichips25_sap3/_1301_ ;
 wire \heichips25_sap3/_1302_ ;
 wire \heichips25_sap3/_1303_ ;
 wire \heichips25_sap3/_1304_ ;
 wire \heichips25_sap3/_1305_ ;
 wire \heichips25_sap3/_1306_ ;
 wire \heichips25_sap3/_1307_ ;
 wire \heichips25_sap3/_1308_ ;
 wire \heichips25_sap3/_1309_ ;
 wire \heichips25_sap3/_1310_ ;
 wire \heichips25_sap3/_1311_ ;
 wire \heichips25_sap3/_1312_ ;
 wire \heichips25_sap3/_1313_ ;
 wire \heichips25_sap3/_1314_ ;
 wire \heichips25_sap3/_1315_ ;
 wire \heichips25_sap3/_1316_ ;
 wire \heichips25_sap3/_1317_ ;
 wire \heichips25_sap3/_1318_ ;
 wire \heichips25_sap3/_1319_ ;
 wire \heichips25_sap3/_1320_ ;
 wire \heichips25_sap3/_1321_ ;
 wire \heichips25_sap3/_1322_ ;
 wire \heichips25_sap3/_1323_ ;
 wire \heichips25_sap3/_1324_ ;
 wire \heichips25_sap3/_1325_ ;
 wire \heichips25_sap3/_1326_ ;
 wire \heichips25_sap3/_1327_ ;
 wire \heichips25_sap3/_1328_ ;
 wire \heichips25_sap3/_1329_ ;
 wire \heichips25_sap3/_1330_ ;
 wire \heichips25_sap3/_1331_ ;
 wire \heichips25_sap3/_1332_ ;
 wire \heichips25_sap3/_1333_ ;
 wire \heichips25_sap3/_1334_ ;
 wire \heichips25_sap3/_1335_ ;
 wire \heichips25_sap3/_1336_ ;
 wire \heichips25_sap3/_1337_ ;
 wire \heichips25_sap3/_1338_ ;
 wire \heichips25_sap3/_1339_ ;
 wire \heichips25_sap3/_1340_ ;
 wire \heichips25_sap3/_1341_ ;
 wire \heichips25_sap3/_1342_ ;
 wire \heichips25_sap3/_1343_ ;
 wire \heichips25_sap3/_1344_ ;
 wire \heichips25_sap3/_1345_ ;
 wire \heichips25_sap3/_1346_ ;
 wire \heichips25_sap3/_1347_ ;
 wire \heichips25_sap3/_1348_ ;
 wire \heichips25_sap3/_1349_ ;
 wire \heichips25_sap3/_1350_ ;
 wire \heichips25_sap3/_1351_ ;
 wire \heichips25_sap3/_1352_ ;
 wire \heichips25_sap3/_1353_ ;
 wire \heichips25_sap3/_1354_ ;
 wire \heichips25_sap3/_1355_ ;
 wire \heichips25_sap3/_1356_ ;
 wire \heichips25_sap3/_1357_ ;
 wire \heichips25_sap3/_1358_ ;
 wire \heichips25_sap3/_1359_ ;
 wire \heichips25_sap3/_1360_ ;
 wire \heichips25_sap3/_1361_ ;
 wire \heichips25_sap3/_1362_ ;
 wire \heichips25_sap3/_1363_ ;
 wire \heichips25_sap3/_1364_ ;
 wire \heichips25_sap3/_1365_ ;
 wire \heichips25_sap3/_1366_ ;
 wire \heichips25_sap3/_1367_ ;
 wire \heichips25_sap3/_1368_ ;
 wire \heichips25_sap3/_1369_ ;
 wire \heichips25_sap3/_1370_ ;
 wire \heichips25_sap3/_1371_ ;
 wire \heichips25_sap3/_1372_ ;
 wire \heichips25_sap3/_1373_ ;
 wire \heichips25_sap3/_1374_ ;
 wire \heichips25_sap3/_1375_ ;
 wire \heichips25_sap3/_1376_ ;
 wire \heichips25_sap3/_1377_ ;
 wire \heichips25_sap3/_1378_ ;
 wire \heichips25_sap3/_1379_ ;
 wire \heichips25_sap3/_1380_ ;
 wire \heichips25_sap3/_1381_ ;
 wire \heichips25_sap3/_1382_ ;
 wire \heichips25_sap3/_1383_ ;
 wire \heichips25_sap3/_1384_ ;
 wire \heichips25_sap3/_1385_ ;
 wire \heichips25_sap3/_1386_ ;
 wire \heichips25_sap3/_1387_ ;
 wire \heichips25_sap3/_1388_ ;
 wire \heichips25_sap3/_1389_ ;
 wire \heichips25_sap3/_1390_ ;
 wire \heichips25_sap3/_1391_ ;
 wire \heichips25_sap3/_1392_ ;
 wire \heichips25_sap3/_1393_ ;
 wire \heichips25_sap3/_1394_ ;
 wire \heichips25_sap3/_1395_ ;
 wire \heichips25_sap3/_1396_ ;
 wire \heichips25_sap3/_1397_ ;
 wire \heichips25_sap3/_1398_ ;
 wire \heichips25_sap3/_1399_ ;
 wire \heichips25_sap3/_1400_ ;
 wire \heichips25_sap3/_1401_ ;
 wire \heichips25_sap3/_1402_ ;
 wire \heichips25_sap3/_1403_ ;
 wire \heichips25_sap3/_1404_ ;
 wire \heichips25_sap3/_1405_ ;
 wire \heichips25_sap3/_1406_ ;
 wire \heichips25_sap3/_1407_ ;
 wire \heichips25_sap3/_1408_ ;
 wire \heichips25_sap3/_1409_ ;
 wire \heichips25_sap3/_1410_ ;
 wire \heichips25_sap3/_1411_ ;
 wire \heichips25_sap3/_1412_ ;
 wire \heichips25_sap3/_1413_ ;
 wire \heichips25_sap3/_1414_ ;
 wire \heichips25_sap3/_1415_ ;
 wire \heichips25_sap3/_1416_ ;
 wire \heichips25_sap3/_1417_ ;
 wire \heichips25_sap3/_1418_ ;
 wire \heichips25_sap3/_1419_ ;
 wire \heichips25_sap3/_1420_ ;
 wire \heichips25_sap3/_1421_ ;
 wire \heichips25_sap3/_1422_ ;
 wire \heichips25_sap3/_1423_ ;
 wire \heichips25_sap3/_1424_ ;
 wire \heichips25_sap3/_1425_ ;
 wire \heichips25_sap3/_1426_ ;
 wire \heichips25_sap3/_1427_ ;
 wire \heichips25_sap3/_1428_ ;
 wire \heichips25_sap3/_1429_ ;
 wire \heichips25_sap3/_1430_ ;
 wire \heichips25_sap3/_1431_ ;
 wire \heichips25_sap3/_1432_ ;
 wire \heichips25_sap3/_1433_ ;
 wire \heichips25_sap3/_1434_ ;
 wire \heichips25_sap3/_1435_ ;
 wire \heichips25_sap3/_1436_ ;
 wire \heichips25_sap3/_1437_ ;
 wire \heichips25_sap3/_1438_ ;
 wire \heichips25_sap3/_1439_ ;
 wire \heichips25_sap3/_1440_ ;
 wire \heichips25_sap3/_1441_ ;
 wire \heichips25_sap3/_1442_ ;
 wire \heichips25_sap3/_1443_ ;
 wire \heichips25_sap3/_1444_ ;
 wire \heichips25_sap3/_1445_ ;
 wire \heichips25_sap3/_1446_ ;
 wire \heichips25_sap3/_1447_ ;
 wire \heichips25_sap3/_1448_ ;
 wire \heichips25_sap3/_1449_ ;
 wire \heichips25_sap3/_1450_ ;
 wire \heichips25_sap3/_1451_ ;
 wire \heichips25_sap3/_1452_ ;
 wire \heichips25_sap3/_1453_ ;
 wire \heichips25_sap3/_1454_ ;
 wire \heichips25_sap3/_1455_ ;
 wire \heichips25_sap3/_1456_ ;
 wire \heichips25_sap3/_1457_ ;
 wire \heichips25_sap3/_1458_ ;
 wire \heichips25_sap3/_1459_ ;
 wire \heichips25_sap3/_1460_ ;
 wire \heichips25_sap3/_1461_ ;
 wire \heichips25_sap3/_1462_ ;
 wire \heichips25_sap3/_1463_ ;
 wire \heichips25_sap3/_1464_ ;
 wire \heichips25_sap3/_1465_ ;
 wire \heichips25_sap3/_1466_ ;
 wire \heichips25_sap3/_1467_ ;
 wire \heichips25_sap3/_1468_ ;
 wire \heichips25_sap3/_1469_ ;
 wire \heichips25_sap3/_1470_ ;
 wire \heichips25_sap3/_1471_ ;
 wire \heichips25_sap3/_1472_ ;
 wire \heichips25_sap3/_1473_ ;
 wire \heichips25_sap3/_1474_ ;
 wire \heichips25_sap3/_1475_ ;
 wire \heichips25_sap3/_1476_ ;
 wire \heichips25_sap3/_1477_ ;
 wire \heichips25_sap3/_1478_ ;
 wire \heichips25_sap3/_1479_ ;
 wire \heichips25_sap3/_1480_ ;
 wire \heichips25_sap3/_1481_ ;
 wire \heichips25_sap3/_1482_ ;
 wire \heichips25_sap3/_1483_ ;
 wire \heichips25_sap3/_1484_ ;
 wire \heichips25_sap3/_1485_ ;
 wire \heichips25_sap3/_1486_ ;
 wire \heichips25_sap3/_1487_ ;
 wire \heichips25_sap3/_1488_ ;
 wire \heichips25_sap3/_1489_ ;
 wire \heichips25_sap3/_1490_ ;
 wire \heichips25_sap3/_1491_ ;
 wire \heichips25_sap3/_1492_ ;
 wire \heichips25_sap3/_1493_ ;
 wire \heichips25_sap3/_1494_ ;
 wire \heichips25_sap3/_1495_ ;
 wire \heichips25_sap3/_1496_ ;
 wire \heichips25_sap3/_1497_ ;
 wire \heichips25_sap3/_1498_ ;
 wire \heichips25_sap3/_1499_ ;
 wire \heichips25_sap3/_1500_ ;
 wire \heichips25_sap3/_1501_ ;
 wire \heichips25_sap3/_1502_ ;
 wire \heichips25_sap3/_1503_ ;
 wire \heichips25_sap3/_1504_ ;
 wire \heichips25_sap3/_1505_ ;
 wire \heichips25_sap3/_1506_ ;
 wire \heichips25_sap3/_1507_ ;
 wire \heichips25_sap3/_1508_ ;
 wire \heichips25_sap3/_1509_ ;
 wire \heichips25_sap3/_1510_ ;
 wire \heichips25_sap3/_1511_ ;
 wire \heichips25_sap3/_1512_ ;
 wire \heichips25_sap3/_1513_ ;
 wire \heichips25_sap3/_1514_ ;
 wire \heichips25_sap3/_1515_ ;
 wire \heichips25_sap3/_1516_ ;
 wire \heichips25_sap3/_1517_ ;
 wire \heichips25_sap3/_1518_ ;
 wire \heichips25_sap3/_1519_ ;
 wire \heichips25_sap3/_1520_ ;
 wire \heichips25_sap3/_1521_ ;
 wire \heichips25_sap3/_1522_ ;
 wire \heichips25_sap3/_1523_ ;
 wire \heichips25_sap3/_1524_ ;
 wire \heichips25_sap3/_1525_ ;
 wire \heichips25_sap3/_1526_ ;
 wire \heichips25_sap3/_1527_ ;
 wire \heichips25_sap3/_1528_ ;
 wire \heichips25_sap3/_1529_ ;
 wire \heichips25_sap3/_1530_ ;
 wire \heichips25_sap3/_1531_ ;
 wire \heichips25_sap3/_1532_ ;
 wire \heichips25_sap3/_1533_ ;
 wire \heichips25_sap3/_1534_ ;
 wire \heichips25_sap3/_1535_ ;
 wire \heichips25_sap3/_1536_ ;
 wire \heichips25_sap3/_1537_ ;
 wire \heichips25_sap3/_1538_ ;
 wire \heichips25_sap3/_1539_ ;
 wire \heichips25_sap3/_1540_ ;
 wire \heichips25_sap3/_1541_ ;
 wire \heichips25_sap3/_1542_ ;
 wire \heichips25_sap3/_1543_ ;
 wire \heichips25_sap3/_1544_ ;
 wire \heichips25_sap3/_1545_ ;
 wire \heichips25_sap3/_1546_ ;
 wire \heichips25_sap3/_1547_ ;
 wire \heichips25_sap3/_1548_ ;
 wire \heichips25_sap3/_1549_ ;
 wire \heichips25_sap3/_1550_ ;
 wire \heichips25_sap3/_1551_ ;
 wire \heichips25_sap3/_1552_ ;
 wire \heichips25_sap3/_1553_ ;
 wire \heichips25_sap3/_1554_ ;
 wire \heichips25_sap3/_1555_ ;
 wire \heichips25_sap3/_1556_ ;
 wire \heichips25_sap3/_1557_ ;
 wire \heichips25_sap3/_1558_ ;
 wire \heichips25_sap3/_1559_ ;
 wire \heichips25_sap3/_1560_ ;
 wire \heichips25_sap3/_1561_ ;
 wire \heichips25_sap3/_1562_ ;
 wire \heichips25_sap3/_1563_ ;
 wire \heichips25_sap3/_1564_ ;
 wire \heichips25_sap3/_1565_ ;
 wire \heichips25_sap3/_1566_ ;
 wire \heichips25_sap3/_1567_ ;
 wire \heichips25_sap3/_1568_ ;
 wire \heichips25_sap3/_1569_ ;
 wire \heichips25_sap3/_1570_ ;
 wire \heichips25_sap3/_1571_ ;
 wire \heichips25_sap3/_1572_ ;
 wire \heichips25_sap3/_1573_ ;
 wire \heichips25_sap3/_1574_ ;
 wire \heichips25_sap3/_1575_ ;
 wire \heichips25_sap3/_1576_ ;
 wire \heichips25_sap3/_1577_ ;
 wire \heichips25_sap3/_1578_ ;
 wire \heichips25_sap3/_1579_ ;
 wire \heichips25_sap3/_1580_ ;
 wire \heichips25_sap3/_1581_ ;
 wire \heichips25_sap3/_1582_ ;
 wire \heichips25_sap3/_1583_ ;
 wire \heichips25_sap3/_1584_ ;
 wire \heichips25_sap3/_1585_ ;
 wire \heichips25_sap3/_1586_ ;
 wire \heichips25_sap3/_1587_ ;
 wire \heichips25_sap3/_1588_ ;
 wire \heichips25_sap3/_1589_ ;
 wire \heichips25_sap3/_1590_ ;
 wire \heichips25_sap3/_1591_ ;
 wire \heichips25_sap3/_1592_ ;
 wire \heichips25_sap3/_1593_ ;
 wire \heichips25_sap3/_1594_ ;
 wire \heichips25_sap3/_1595_ ;
 wire \heichips25_sap3/_1596_ ;
 wire \heichips25_sap3/_1597_ ;
 wire \heichips25_sap3/_1598_ ;
 wire \heichips25_sap3/_1599_ ;
 wire \heichips25_sap3/_1600_ ;
 wire \heichips25_sap3/_1601_ ;
 wire \heichips25_sap3/_1602_ ;
 wire \heichips25_sap3/_1603_ ;
 wire \heichips25_sap3/_1604_ ;
 wire \heichips25_sap3/_1605_ ;
 wire \heichips25_sap3/_1606_ ;
 wire \heichips25_sap3/_1607_ ;
 wire \heichips25_sap3/_1608_ ;
 wire \heichips25_sap3/_1609_ ;
 wire \heichips25_sap3/_1610_ ;
 wire \heichips25_sap3/_1611_ ;
 wire \heichips25_sap3/_1612_ ;
 wire \heichips25_sap3/_1613_ ;
 wire \heichips25_sap3/_1614_ ;
 wire \heichips25_sap3/_1615_ ;
 wire \heichips25_sap3/_1616_ ;
 wire \heichips25_sap3/_1617_ ;
 wire \heichips25_sap3/_1618_ ;
 wire \heichips25_sap3/_1619_ ;
 wire \heichips25_sap3/_1620_ ;
 wire \heichips25_sap3/_1621_ ;
 wire \heichips25_sap3/_1622_ ;
 wire \heichips25_sap3/_1623_ ;
 wire \heichips25_sap3/_1624_ ;
 wire \heichips25_sap3/_1625_ ;
 wire \heichips25_sap3/_1626_ ;
 wire \heichips25_sap3/_1627_ ;
 wire \heichips25_sap3/_1628_ ;
 wire \heichips25_sap3/_1629_ ;
 wire \heichips25_sap3/_1630_ ;
 wire \heichips25_sap3/_1631_ ;
 wire \heichips25_sap3/_1632_ ;
 wire \heichips25_sap3/_1633_ ;
 wire \heichips25_sap3/_1634_ ;
 wire \heichips25_sap3/_1635_ ;
 wire \heichips25_sap3/_1636_ ;
 wire \heichips25_sap3/_1637_ ;
 wire \heichips25_sap3/_1638_ ;
 wire \heichips25_sap3/_1639_ ;
 wire \heichips25_sap3/_1640_ ;
 wire \heichips25_sap3/_1641_ ;
 wire \heichips25_sap3/_1642_ ;
 wire \heichips25_sap3/_1643_ ;
 wire \heichips25_sap3/_1644_ ;
 wire \heichips25_sap3/_1645_ ;
 wire \heichips25_sap3/_1646_ ;
 wire \heichips25_sap3/_1647_ ;
 wire \heichips25_sap3/_1648_ ;
 wire \heichips25_sap3/_1649_ ;
 wire \heichips25_sap3/_1650_ ;
 wire \heichips25_sap3/_1651_ ;
 wire \heichips25_sap3/_1652_ ;
 wire \heichips25_sap3/_1653_ ;
 wire \heichips25_sap3/_1654_ ;
 wire \heichips25_sap3/_1655_ ;
 wire \heichips25_sap3/_1656_ ;
 wire \heichips25_sap3/_1657_ ;
 wire \heichips25_sap3/_1658_ ;
 wire \heichips25_sap3/_1659_ ;
 wire \heichips25_sap3/_1660_ ;
 wire \heichips25_sap3/_1661_ ;
 wire \heichips25_sap3/_1662_ ;
 wire \heichips25_sap3/_1663_ ;
 wire \heichips25_sap3/_1664_ ;
 wire \heichips25_sap3/_1665_ ;
 wire \heichips25_sap3/_1666_ ;
 wire \heichips25_sap3/_1667_ ;
 wire \heichips25_sap3/_1668_ ;
 wire \heichips25_sap3/_1669_ ;
 wire \heichips25_sap3/_1670_ ;
 wire \heichips25_sap3/_1671_ ;
 wire \heichips25_sap3/_1672_ ;
 wire \heichips25_sap3/_1673_ ;
 wire \heichips25_sap3/_1674_ ;
 wire \heichips25_sap3/_1675_ ;
 wire \heichips25_sap3/_1676_ ;
 wire \heichips25_sap3/_1677_ ;
 wire \heichips25_sap3/_1678_ ;
 wire \heichips25_sap3/_1679_ ;
 wire \heichips25_sap3/_1680_ ;
 wire \heichips25_sap3/_1681_ ;
 wire \heichips25_sap3/_1682_ ;
 wire \heichips25_sap3/_1683_ ;
 wire \heichips25_sap3/_1684_ ;
 wire \heichips25_sap3/_1685_ ;
 wire \heichips25_sap3/_1686_ ;
 wire \heichips25_sap3/_1687_ ;
 wire \heichips25_sap3/_1688_ ;
 wire \heichips25_sap3/_1689_ ;
 wire \heichips25_sap3/_1690_ ;
 wire \heichips25_sap3/_1691_ ;
 wire \heichips25_sap3/_1692_ ;
 wire \heichips25_sap3/_1693_ ;
 wire \heichips25_sap3/_1694_ ;
 wire \heichips25_sap3/_1695_ ;
 wire \heichips25_sap3/_1696_ ;
 wire \heichips25_sap3/_1697_ ;
 wire \heichips25_sap3/_1698_ ;
 wire \heichips25_sap3/_1699_ ;
 wire \heichips25_sap3/_1700_ ;
 wire \heichips25_sap3/_1701_ ;
 wire \heichips25_sap3/_1702_ ;
 wire \heichips25_sap3/_1703_ ;
 wire \heichips25_sap3/_1704_ ;
 wire \heichips25_sap3/_1705_ ;
 wire \heichips25_sap3/_1706_ ;
 wire \heichips25_sap3/_1707_ ;
 wire \heichips25_sap3/_1708_ ;
 wire \heichips25_sap3/_1709_ ;
 wire \heichips25_sap3/_1710_ ;
 wire \heichips25_sap3/_1711_ ;
 wire \heichips25_sap3/_1712_ ;
 wire \heichips25_sap3/_1713_ ;
 wire \heichips25_sap3/_1714_ ;
 wire \heichips25_sap3/_1715_ ;
 wire \heichips25_sap3/_1716_ ;
 wire \heichips25_sap3/_1717_ ;
 wire \heichips25_sap3/_1718_ ;
 wire \heichips25_sap3/_1719_ ;
 wire \heichips25_sap3/_1720_ ;
 wire \heichips25_sap3/_1721_ ;
 wire \heichips25_sap3/_1722_ ;
 wire \heichips25_sap3/_1723_ ;
 wire \heichips25_sap3/_1724_ ;
 wire \heichips25_sap3/_1725_ ;
 wire \heichips25_sap3/_1726_ ;
 wire \heichips25_sap3/_1727_ ;
 wire \heichips25_sap3/_1728_ ;
 wire \heichips25_sap3/_1729_ ;
 wire \heichips25_sap3/_1730_ ;
 wire \heichips25_sap3/_1731_ ;
 wire \heichips25_sap3/_1732_ ;
 wire \heichips25_sap3/_1733_ ;
 wire \heichips25_sap3/_1734_ ;
 wire \heichips25_sap3/_1735_ ;
 wire \heichips25_sap3/_1736_ ;
 wire \heichips25_sap3/_1737_ ;
 wire \heichips25_sap3/_1738_ ;
 wire \heichips25_sap3/_1739_ ;
 wire \heichips25_sap3/_1740_ ;
 wire \heichips25_sap3/_1741_ ;
 wire \heichips25_sap3/_1742_ ;
 wire \heichips25_sap3/_1743_ ;
 wire \heichips25_sap3/_1744_ ;
 wire \heichips25_sap3/_1745_ ;
 wire \heichips25_sap3/_1746_ ;
 wire \heichips25_sap3/_1747_ ;
 wire \heichips25_sap3/_1748_ ;
 wire \heichips25_sap3/_1749_ ;
 wire \heichips25_sap3/_1750_ ;
 wire \heichips25_sap3/_1751_ ;
 wire \heichips25_sap3/_1752_ ;
 wire \heichips25_sap3/_1753_ ;
 wire \heichips25_sap3/_1754_ ;
 wire \heichips25_sap3/_1755_ ;
 wire \heichips25_sap3/_1756_ ;
 wire \heichips25_sap3/_1757_ ;
 wire \heichips25_sap3/_1758_ ;
 wire \heichips25_sap3/_1759_ ;
 wire \heichips25_sap3/_1760_ ;
 wire \heichips25_sap3/_1761_ ;
 wire \heichips25_sap3/_1762_ ;
 wire \heichips25_sap3/_1763_ ;
 wire \heichips25_sap3/_1764_ ;
 wire \heichips25_sap3/_1765_ ;
 wire \heichips25_sap3/_1766_ ;
 wire \heichips25_sap3/_1767_ ;
 wire \heichips25_sap3/_1768_ ;
 wire \heichips25_sap3/_1769_ ;
 wire \heichips25_sap3/_1770_ ;
 wire \heichips25_sap3/_1771_ ;
 wire \heichips25_sap3/_1772_ ;
 wire \heichips25_sap3/_1773_ ;
 wire \heichips25_sap3/_1774_ ;
 wire \heichips25_sap3/_1775_ ;
 wire \heichips25_sap3/_1776_ ;
 wire \heichips25_sap3/_1777_ ;
 wire \heichips25_sap3/_1778_ ;
 wire \heichips25_sap3/_1779_ ;
 wire \heichips25_sap3/_1780_ ;
 wire \heichips25_sap3/_1781_ ;
 wire \heichips25_sap3/_1782_ ;
 wire \heichips25_sap3/_1783_ ;
 wire \heichips25_sap3/_1784_ ;
 wire \heichips25_sap3/_1785_ ;
 wire \heichips25_sap3/_1786_ ;
 wire \heichips25_sap3/_1787_ ;
 wire \heichips25_sap3/_1788_ ;
 wire \heichips25_sap3/_1789_ ;
 wire \heichips25_sap3/_1790_ ;
 wire \heichips25_sap3/_1791_ ;
 wire \heichips25_sap3/_1792_ ;
 wire \heichips25_sap3/_1793_ ;
 wire \heichips25_sap3/_1794_ ;
 wire \heichips25_sap3/_1795_ ;
 wire \heichips25_sap3/_1796_ ;
 wire \heichips25_sap3/_1797_ ;
 wire \heichips25_sap3/_1798_ ;
 wire \heichips25_sap3/_1799_ ;
 wire \heichips25_sap3/_1800_ ;
 wire \heichips25_sap3/_1801_ ;
 wire \heichips25_sap3/_1802_ ;
 wire \heichips25_sap3/_1803_ ;
 wire \heichips25_sap3/_1804_ ;
 wire \heichips25_sap3/_1805_ ;
 wire \heichips25_sap3/_1806_ ;
 wire \heichips25_sap3/_1807_ ;
 wire \heichips25_sap3/_1808_ ;
 wire \heichips25_sap3/_1809_ ;
 wire \heichips25_sap3/_1810_ ;
 wire \heichips25_sap3/_1811_ ;
 wire \heichips25_sap3/_1812_ ;
 wire \heichips25_sap3/_1813_ ;
 wire \heichips25_sap3/_1814_ ;
 wire \heichips25_sap3/_1815_ ;
 wire \heichips25_sap3/_1816_ ;
 wire \heichips25_sap3/_1817_ ;
 wire \heichips25_sap3/_1818_ ;
 wire \heichips25_sap3/_1819_ ;
 wire \heichips25_sap3/_1820_ ;
 wire \heichips25_sap3/_1821_ ;
 wire \heichips25_sap3/_1822_ ;
 wire \heichips25_sap3/_1823_ ;
 wire \heichips25_sap3/_1824_ ;
 wire \heichips25_sap3/_1825_ ;
 wire \heichips25_sap3/_1826_ ;
 wire \heichips25_sap3/_1827_ ;
 wire \heichips25_sap3/_1828_ ;
 wire \heichips25_sap3/_1829_ ;
 wire \heichips25_sap3/_1830_ ;
 wire \heichips25_sap3/_1831_ ;
 wire \heichips25_sap3/_1832_ ;
 wire \heichips25_sap3/_1833_ ;
 wire \heichips25_sap3/_1834_ ;
 wire \heichips25_sap3/_1835_ ;
 wire \heichips25_sap3/_1836_ ;
 wire \heichips25_sap3/_1837_ ;
 wire \heichips25_sap3/_1838_ ;
 wire \heichips25_sap3/_1839_ ;
 wire \heichips25_sap3/_1840_ ;
 wire \heichips25_sap3/_1841_ ;
 wire \heichips25_sap3/_1842_ ;
 wire \heichips25_sap3/_1843_ ;
 wire \heichips25_sap3/_1844_ ;
 wire \heichips25_sap3/_1845_ ;
 wire \heichips25_sap3/_1846_ ;
 wire \heichips25_sap3/_1847_ ;
 wire \heichips25_sap3/_1848_ ;
 wire \heichips25_sap3/_1849_ ;
 wire \heichips25_sap3/_1850_ ;
 wire \heichips25_sap3/_1851_ ;
 wire \heichips25_sap3/_1852_ ;
 wire \heichips25_sap3/_1853_ ;
 wire \heichips25_sap3/_1854_ ;
 wire \heichips25_sap3/_1855_ ;
 wire \heichips25_sap3/_1856_ ;
 wire \heichips25_sap3/_1857_ ;
 wire \heichips25_sap3/_1858_ ;
 wire \heichips25_sap3/_1859_ ;
 wire \heichips25_sap3/_1860_ ;
 wire \heichips25_sap3/_1861_ ;
 wire \heichips25_sap3/_1862_ ;
 wire \heichips25_sap3/_1863_ ;
 wire \heichips25_sap3/_1864_ ;
 wire \heichips25_sap3/_1865_ ;
 wire \heichips25_sap3/_1866_ ;
 wire \heichips25_sap3/_1867_ ;
 wire \heichips25_sap3/_1868_ ;
 wire \heichips25_sap3/_1869_ ;
 wire \heichips25_sap3/_1870_ ;
 wire \heichips25_sap3/_1871_ ;
 wire \heichips25_sap3/_1872_ ;
 wire \heichips25_sap3/_1873_ ;
 wire \heichips25_sap3/_1874_ ;
 wire \heichips25_sap3/_1875_ ;
 wire \heichips25_sap3/_1876_ ;
 wire \heichips25_sap3/_1877_ ;
 wire \heichips25_sap3/_1878_ ;
 wire \heichips25_sap3/_1879_ ;
 wire \heichips25_sap3/_1880_ ;
 wire \heichips25_sap3/_1881_ ;
 wire \heichips25_sap3/_1882_ ;
 wire \heichips25_sap3/_1883_ ;
 wire \heichips25_sap3/_1884_ ;
 wire \heichips25_sap3/_1885_ ;
 wire \heichips25_sap3/_1886_ ;
 wire \heichips25_sap3/_1887_ ;
 wire \heichips25_sap3/_1888_ ;
 wire \heichips25_sap3/_1889_ ;
 wire \heichips25_sap3/_1890_ ;
 wire \heichips25_sap3/_1891_ ;
 wire \heichips25_sap3/_1892_ ;
 wire \heichips25_sap3/_1893_ ;
 wire \heichips25_sap3/_1894_ ;
 wire \heichips25_sap3/_1895_ ;
 wire \heichips25_sap3/_1896_ ;
 wire \heichips25_sap3/_1897_ ;
 wire \heichips25_sap3/_1898_ ;
 wire \heichips25_sap3/_1899_ ;
 wire \heichips25_sap3/_1900_ ;
 wire \heichips25_sap3/_1901_ ;
 wire \heichips25_sap3/_1902_ ;
 wire \heichips25_sap3/_1903_ ;
 wire \heichips25_sap3/_1904_ ;
 wire \heichips25_sap3/_1905_ ;
 wire \heichips25_sap3/_1906_ ;
 wire \heichips25_sap3/_1907_ ;
 wire \heichips25_sap3/_1908_ ;
 wire \heichips25_sap3/_1909_ ;
 wire \heichips25_sap3/_1910_ ;
 wire \heichips25_sap3/_1911_ ;
 wire \heichips25_sap3/_1912_ ;
 wire \heichips25_sap3/_1913_ ;
 wire \heichips25_sap3/_1914_ ;
 wire \heichips25_sap3/_1915_ ;
 wire \heichips25_sap3/_1916_ ;
 wire \heichips25_sap3/_1917_ ;
 wire \heichips25_sap3/_1918_ ;
 wire \heichips25_sap3/_1919_ ;
 wire \heichips25_sap3/_1920_ ;
 wire \heichips25_sap3/_1921_ ;
 wire \heichips25_sap3/_1922_ ;
 wire \heichips25_sap3/_1923_ ;
 wire \heichips25_sap3/_1924_ ;
 wire \heichips25_sap3/_1925_ ;
 wire \heichips25_sap3/_1926_ ;
 wire \heichips25_sap3/_1927_ ;
 wire \heichips25_sap3/_1928_ ;
 wire \heichips25_sap3/_1929_ ;
 wire \heichips25_sap3/_1930_ ;
 wire \heichips25_sap3/_1931_ ;
 wire \heichips25_sap3/clk_div_out ;
 wire \heichips25_sap3/mem_mar_we ;
 wire \heichips25_sap3/mem_ram_we ;
 wire \heichips25_sap3/regFile_serial ;
 wire \heichips25_sap3/regFile_serial_start ;
 wire \heichips25_sap3/sap_3_inst.alu_flags[0] ;
 wire \heichips25_sap3/sap_3_inst.alu_flags[1] ;
 wire \heichips25_sap3/sap_3_inst.alu_flags[2] ;
 wire \heichips25_sap3/sap_3_inst.alu_flags[3] ;
 wire \heichips25_sap3/sap_3_inst.alu_flags[4] ;
 wire \heichips25_sap3/sap_3_inst.alu_flags[5] ;
 wire \heichips25_sap3/sap_3_inst.alu_flags[6] ;
 wire \heichips25_sap3/sap_3_inst.alu_flags[7] ;
 wire \heichips25_sap3/sap_3_inst.alu_inst.acc[0] ;
 wire \heichips25_sap3/sap_3_inst.alu_inst.acc[1] ;
 wire \heichips25_sap3/sap_3_inst.alu_inst.acc[2] ;
 wire \heichips25_sap3/sap_3_inst.alu_inst.acc[3] ;
 wire \heichips25_sap3/sap_3_inst.alu_inst.acc[4] ;
 wire \heichips25_sap3/sap_3_inst.alu_inst.acc[5] ;
 wire \heichips25_sap3/sap_3_inst.alu_inst.acc[6] ;
 wire \heichips25_sap3/sap_3_inst.alu_inst.acc[7] ;
 wire \heichips25_sap3/sap_3_inst.alu_inst.act[0] ;
 wire \heichips25_sap3/sap_3_inst.alu_inst.act[1] ;
 wire \heichips25_sap3/sap_3_inst.alu_inst.act[2] ;
 wire \heichips25_sap3/sap_3_inst.alu_inst.act[3] ;
 wire \heichips25_sap3/sap_3_inst.alu_inst.act[4] ;
 wire \heichips25_sap3/sap_3_inst.alu_inst.act[5] ;
 wire \heichips25_sap3/sap_3_inst.alu_inst.act[6] ;
 wire \heichips25_sap3/sap_3_inst.alu_inst.act[7] ;
 wire \heichips25_sap3/sap_3_inst.alu_inst.carry ;
 wire \heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \heichips25_sap3/sap_3_inst.alu_inst.tmp[0] ;
 wire \heichips25_sap3/sap_3_inst.alu_inst.tmp[1] ;
 wire \heichips25_sap3/sap_3_inst.alu_inst.tmp[2] ;
 wire \heichips25_sap3/sap_3_inst.alu_inst.tmp[3] ;
 wire \heichips25_sap3/sap_3_inst.alu_inst.tmp[4] ;
 wire \heichips25_sap3/sap_3_inst.alu_inst.tmp[5] ;
 wire \heichips25_sap3/sap_3_inst.alu_inst.tmp[6] ;
 wire \heichips25_sap3/sap_3_inst.alu_inst.tmp[7] ;
 wire \heichips25_sap3/sap_3_inst.controller_inst.opcode[0] ;
 wire \heichips25_sap3/sap_3_inst.controller_inst.opcode[1] ;
 wire \heichips25_sap3/sap_3_inst.controller_inst.opcode[2] ;
 wire \heichips25_sap3/sap_3_inst.controller_inst.opcode[3] ;
 wire \heichips25_sap3/sap_3_inst.controller_inst.opcode[4] ;
 wire \heichips25_sap3/sap_3_inst.controller_inst.opcode[5] ;
 wire \heichips25_sap3/sap_3_inst.controller_inst.opcode[6] ;
 wire \heichips25_sap3/sap_3_inst.controller_inst.opcode[7] ;
 wire \heichips25_sap3/sap_3_inst.controller_inst.stage[0] ;
 wire \heichips25_sap3/sap_3_inst.controller_inst.stage[1] ;
 wire \heichips25_sap3/sap_3_inst.controller_inst.stage[2] ;
 wire \heichips25_sap3/sap_3_inst.controller_inst.stage[3] ;
 wire \heichips25_sap3/sap_3_inst.out[0] ;
 wire \heichips25_sap3/sap_3_inst.out[1] ;
 wire \heichips25_sap3/sap_3_inst.out[2] ;
 wire \heichips25_sap3/sap_3_inst.out[3] ;
 wire \heichips25_sap3/sap_3_inst.out[4] ;
 wire \heichips25_sap3/sap_3_inst.out[5] ;
 wire \heichips25_sap3/sap_3_inst.out[6] ;
 wire \heichips25_sap3/sap_3_inst.out[7] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos[0] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos[1] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos[2] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[0][0] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[0][1] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[0][2] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[0][3] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[0][4] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[0][5] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[0][6] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[0][7] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][0] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][1] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][2] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][3] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][4] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][5] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][6] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][7] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][0] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][1] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][2] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][3] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][4] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][5] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][6] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][7] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][0] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][1] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][2] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][3] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][4] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][5] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][6] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][7] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][0] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][1] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][2] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][3] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][4] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][5] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][6] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][7] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][0] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][1] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][2] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][3] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][4] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][5] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][6] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][7] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][0] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][1] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][2] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][3] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][4] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][5] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][6] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][7] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][0] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][1] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][2] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][3] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][4] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][5] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][6] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][7] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][0] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][1] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][2] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][3] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][4] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][5] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][6] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][7] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][0] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][1] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][2] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][3] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][4] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][5] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][6] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][7] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][0] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][1] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][2] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][3] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][4] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][5] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][6] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][7] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][0] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][1] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][2] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][3] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][4] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][5] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][6] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][7] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[0] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[1] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[2] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[3] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[4] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[5] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[6] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[7] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.state[0] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.state[1] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.state[2] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.word_index[0] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.word_index[1] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.word_index[2] ;
 wire \heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.word_index[3] ;
 wire \heichips25_sap3/sap_3_outputReg_serial ;
 wire \heichips25_sap3/sap_3_outputReg_start_sync ;
 wire \heichips25_sap3/u_ser.bit_pos[0] ;
 wire \heichips25_sap3/u_ser.bit_pos[1] ;
 wire \heichips25_sap3/u_ser.bit_pos[2] ;
 wire \heichips25_sap3/u_ser.shadow_reg[0] ;
 wire \heichips25_sap3/u_ser.shadow_reg[1] ;
 wire \heichips25_sap3/u_ser.shadow_reg[2] ;
 wire \heichips25_sap3/u_ser.shadow_reg[3] ;
 wire \heichips25_sap3/u_ser.shadow_reg[4] ;
 wire \heichips25_sap3/u_ser.shadow_reg[5] ;
 wire \heichips25_sap3/u_ser.shadow_reg[6] ;
 wire \heichips25_sap3/u_ser.shadow_reg[7] ;
 wire \heichips25_sap3/u_ser.state[0] ;
 wire \heichips25_sap3/u_ser.state[1] ;
 wire \heichips25_sap3/u_ser.state[2] ;
 wire \heichips25_sap3/clk_div_param_inst/_0_ ;
 wire \heichips25_sap3/clk_div_param_inst/clk_out_reg ;
 wire net43;
 wire net44;
 wire \heichips25_sap3/net45 ;
 wire net46;
 wire net47;
 wire \heichips25_sap3/net48 ;
 wire \heichips25_sap3/net49 ;
 wire \heichips25_sap3/net50 ;
 wire \heichips25_sap3/net51 ;
 wire \heichips25_sap3/net52 ;
 wire \heichips25_sap3/net53 ;
 wire \heichips25_sap3/net54 ;
 wire \heichips25_sap3/net55 ;
 wire \heichips25_sap3/net56 ;
 wire \heichips25_sap3/net57 ;
 wire \heichips25_sap3/net58 ;
 wire \heichips25_sap3/net59 ;
 wire \heichips25_sap3/net60 ;
 wire \heichips25_sap3/net61 ;
 wire \heichips25_sap3/net62 ;
 wire \heichips25_sap3/net63 ;
 wire \heichips25_sap3/net64 ;
 wire \heichips25_sap3/net65 ;
 wire \heichips25_sap3/net66 ;
 wire \heichips25_sap3/net67 ;
 wire \heichips25_sap3/net68 ;
 wire \heichips25_sap3/net69 ;
 wire \heichips25_sap3/net70 ;
 wire \heichips25_sap3/net71 ;
 wire \heichips25_sap3/net72 ;
 wire \heichips25_sap3/net73 ;
 wire \heichips25_sap3/net74 ;
 wire \heichips25_sap3/net75 ;
 wire \heichips25_sap3/net76 ;
 wire \heichips25_sap3/net77 ;
 wire \heichips25_sap3/net78 ;
 wire \heichips25_sap3/net79 ;
 wire \heichips25_sap3/net80 ;
 wire \heichips25_sap3/net81 ;
 wire \heichips25_sap3/net82 ;
 wire \heichips25_sap3/net83 ;
 wire \heichips25_sap3/net84 ;
 wire \heichips25_sap3/net85 ;
 wire \heichips25_sap3/net86 ;
 wire \heichips25_sap3/net87 ;
 wire \heichips25_sap3/net88 ;
 wire \heichips25_sap3/net89 ;
 wire \heichips25_sap3/net90 ;
 wire \heichips25_sap3/net91 ;
 wire \heichips25_sap3/net92 ;
 wire \heichips25_sap3/net93 ;
 wire \heichips25_sap3/net94 ;
 wire \heichips25_sap3/net95 ;
 wire \heichips25_sap3/net96 ;
 wire \heichips25_sap3/net97 ;
 wire \heichips25_sap3/net98 ;
 wire \heichips25_sap3/net99 ;
 wire \heichips25_sap3/net100 ;
 wire \heichips25_sap3/net101 ;
 wire \heichips25_sap3/net102 ;
 wire \heichips25_sap3/net103 ;
 wire \heichips25_sap3/net104 ;
 wire \heichips25_sap3/net105 ;
 wire \heichips25_sap3/net106 ;
 wire \heichips25_sap3/net107 ;
 wire \heichips25_sap3/net108 ;
 wire \heichips25_sap3/net109 ;
 wire \heichips25_sap3/net110 ;
 wire \heichips25_sap3/net111 ;
 wire \heichips25_sap3/net112 ;
 wire \heichips25_sap3/net113 ;
 wire \heichips25_sap3/net114 ;
 wire \heichips25_sap3/net115 ;
 wire \heichips25_sap3/net116 ;
 wire \heichips25_sap3/net117 ;
 wire \heichips25_sap3/net118 ;
 wire \heichips25_sap3/net119 ;
 wire \heichips25_sap3/net120 ;
 wire \heichips25_sap3/net121 ;
 wire \heichips25_sap3/net122 ;
 wire \heichips25_sap3/net123 ;
 wire \heichips25_sap3/net124 ;
 wire \heichips25_sap3/net125 ;
 wire \heichips25_sap3/net126 ;
 wire \heichips25_sap3/net127 ;
 wire \heichips25_sap3/net128 ;
 wire \heichips25_sap3/net129 ;
 wire \heichips25_sap3/net130 ;
 wire \heichips25_sap3/net131 ;
 wire \heichips25_sap3/net132 ;
 wire \heichips25_sap3/net133 ;
 wire \heichips25_sap3/net134 ;
 wire \heichips25_sap3/net135 ;
 wire \heichips25_sap3/net136 ;
 wire \heichips25_sap3/net137 ;
 wire \heichips25_sap3/net138 ;
 wire \heichips25_sap3/net139 ;
 wire \heichips25_sap3/net140 ;
 wire \heichips25_sap3/net141 ;
 wire \heichips25_sap3/net142 ;
 wire \heichips25_sap3/net143 ;
 wire \heichips25_sap3/net144 ;
 wire \heichips25_sap3/net145 ;
 wire \heichips25_sap3/net146 ;
 wire \heichips25_sap3/net147 ;
 wire \heichips25_sap3/net148 ;
 wire \heichips25_sap3/net149 ;
 wire \heichips25_sap3/net150 ;
 wire \heichips25_sap3/net151 ;
 wire \heichips25_sap3/net152 ;
 wire \heichips25_sap3/net153 ;
 wire \heichips25_sap3/net154 ;
 wire \heichips25_sap3/net155 ;
 wire \heichips25_sap3/net156 ;
 wire \heichips25_sap3/net157 ;
 wire \heichips25_sap3/net158 ;
 wire \heichips25_sap3/net159 ;
 wire \heichips25_can_lehmann_fsm/net160 ;
 wire \heichips25_can_lehmann_fsm/net161 ;
 wire \heichips25_can_lehmann_fsm/net162 ;
 wire \heichips25_can_lehmann_fsm/net163 ;
 wire \heichips25_can_lehmann_fsm/net164 ;
 wire \heichips25_can_lehmann_fsm/net165 ;
 wire \heichips25_sap3/net166 ;
 wire \heichips25_sap3/net167 ;
 wire \heichips25_sap3/net168 ;
 wire \heichips25_sap3/net169 ;
 wire \heichips25_can_lehmann_fsm/net170 ;
 wire \heichips25_can_lehmann_fsm/net171 ;
 wire \heichips25_can_lehmann_fsm/net172 ;
 wire \heichips25_can_lehmann_fsm/net173 ;
 wire \heichips25_can_lehmann_fsm/net174 ;
 wire \heichips25_can_lehmann_fsm/net175 ;
 wire \heichips25_can_lehmann_fsm/net176 ;
 wire \heichips25_can_lehmann_fsm/net177 ;
 wire \heichips25_can_lehmann_fsm/net178 ;
 wire \heichips25_can_lehmann_fsm/net179 ;
 wire \heichips25_can_lehmann_fsm/net180 ;
 wire \heichips25_can_lehmann_fsm/net181 ;
 wire \heichips25_can_lehmann_fsm/net182 ;
 wire \heichips25_can_lehmann_fsm/net183 ;
 wire \heichips25_can_lehmann_fsm/net184 ;
 wire \heichips25_can_lehmann_fsm/net185 ;
 wire \heichips25_can_lehmann_fsm/net186 ;
 wire \heichips25_can_lehmann_fsm/net187 ;
 wire \heichips25_can_lehmann_fsm/net188 ;
 wire \heichips25_can_lehmann_fsm/net189 ;
 wire \heichips25_can_lehmann_fsm/net190 ;
 wire \heichips25_can_lehmann_fsm/net191 ;
 wire \heichips25_can_lehmann_fsm/net192 ;
 wire \heichips25_can_lehmann_fsm/net193 ;
 wire \heichips25_can_lehmann_fsm/net194 ;
 wire \heichips25_can_lehmann_fsm/net195 ;
 wire \heichips25_can_lehmann_fsm/net196 ;
 wire \heichips25_can_lehmann_fsm/net197 ;
 wire \heichips25_can_lehmann_fsm/net198 ;
 wire \heichips25_can_lehmann_fsm/net199 ;
 wire \heichips25_can_lehmann_fsm/net200 ;
 wire \heichips25_sap3/net201 ;
 wire \heichips25_sap3/net202 ;
 wire \heichips25_sap3/net203 ;
 wire \heichips25_sap3/net204 ;
 wire \heichips25_can_lehmann_fsm/net205 ;
 wire \heichips25_can_lehmann_fsm/net206 ;
 wire \heichips25_can_lehmann_fsm/net207 ;
 wire \heichips25_can_lehmann_fsm/net208 ;
 wire \heichips25_can_lehmann_fsm/net209 ;
 wire \heichips25_can_lehmann_fsm/net210 ;
 wire \heichips25_sap3/net211 ;
 wire \heichips25_sap3/net212 ;
 wire \heichips25_sap3/net213 ;
 wire \heichips25_sap3/net214 ;
 wire \heichips25_sap3/net215 ;
 wire \heichips25_sap3/net216 ;
 wire \heichips25_sap3/net217 ;
 wire \heichips25_sap3/net218 ;
 wire \heichips25_can_lehmann_fsm/net219 ;
 wire \heichips25_sap3/net220 ;
 wire \heichips25_sap3/net221 ;
 wire \heichips25_sap3/net222 ;
 wire \heichips25_sap3/net223 ;
 wire \heichips25_sap3/net224 ;
 wire \heichips25_sap3/net225 ;
 wire \heichips25_sap3/net226 ;
 wire \heichips25_sap3/net227 ;
 wire \heichips25_sap3/net228 ;
 wire \heichips25_sap3/net229 ;
 wire \heichips25_sap3/net230 ;
 wire \heichips25_sap3/net231 ;
 wire \heichips25_sap3/net232 ;
 wire \heichips25_sap3/net233 ;
 wire \heichips25_sap3/net234 ;
 wire \heichips25_sap3/net235 ;
 wire \heichips25_sap3/net236 ;
 wire \heichips25_sap3/net237 ;
 wire \heichips25_sap3/net238 ;
 wire \heichips25_sap3/net239 ;
 wire \heichips25_sap3/net240 ;
 wire \heichips25_sap3/net241 ;
 wire \heichips25_sap3/net242 ;
 wire \heichips25_sap3/net243 ;
 wire \heichips25_sap3/net244 ;
 wire \heichips25_sap3/net245 ;
 wire \heichips25_sap3/net246 ;
 wire \heichips25_sap3/net247 ;
 wire \heichips25_sap3/net248 ;
 wire \heichips25_sap3/net249 ;
 wire \heichips25_sap3/net250 ;
 wire \heichips25_sap3/net251 ;
 wire \heichips25_sap3/net252 ;
 wire \heichips25_sap3/net253 ;
 wire \heichips25_sap3/net254 ;
 wire \heichips25_sap3/net255 ;
 wire \heichips25_sap3/net256 ;
 wire \heichips25_sap3/net257 ;
 wire \heichips25_sap3/net258 ;
 wire \heichips25_sap3/net259 ;
 wire \heichips25_sap3/net260 ;
 wire \heichips25_sap3/net261 ;
 wire \heichips25_sap3/net262 ;
 wire \heichips25_sap3/net263 ;
 wire \heichips25_sap3/net264 ;
 wire \heichips25_sap3/net265 ;
 wire \heichips25_sap3/net266 ;
 wire \heichips25_sap3/net267 ;
 wire \heichips25_sap3/net268 ;
 wire \heichips25_sap3/net269 ;
 wire \heichips25_sap3/net270 ;
 wire \heichips25_sap3/net271 ;
 wire \heichips25_sap3/net272 ;
 wire \heichips25_sap3/net273 ;
 wire \heichips25_sap3/net274 ;
 wire \heichips25_sap3/net275 ;
 wire \heichips25_sap3/net276 ;
 wire \heichips25_sap3/net277 ;
 wire \heichips25_sap3/net278 ;
 wire \heichips25_sap3/net279 ;
 wire \heichips25_sap3/net280 ;
 wire \heichips25_sap3/net281 ;
 wire \heichips25_sap3/net282 ;
 wire \heichips25_sap3/net283 ;
 wire \heichips25_sap3/net284 ;
 wire \heichips25_sap3/net285 ;
 wire \heichips25_sap3/net286 ;
 wire \heichips25_sap3/net287 ;
 wire \heichips25_sap3/net288 ;
 wire \heichips25_sap3/net289 ;
 wire \heichips25_sap3/net290 ;
 wire \heichips25_sap3/net291 ;
 wire \heichips25_sap3/net292 ;
 wire \heichips25_sap3/net293 ;
 wire \heichips25_can_lehmann_fsm/net294 ;
 wire \heichips25_can_lehmann_fsm/net295 ;
 wire \heichips25_can_lehmann_fsm/net296 ;
 wire \heichips25_can_lehmann_fsm/net297 ;
 wire \heichips25_can_lehmann_fsm/net298 ;
 wire \heichips25_can_lehmann_fsm/net299 ;
 wire \heichips25_can_lehmann_fsm/net300 ;
 wire \heichips25_can_lehmann_fsm/net301 ;
 wire \heichips25_can_lehmann_fsm/net302 ;
 wire \heichips25_can_lehmann_fsm/net303 ;
 wire \heichips25_can_lehmann_fsm/net304 ;
 wire \heichips25_can_lehmann_fsm/net305 ;
 wire \heichips25_can_lehmann_fsm/net306 ;
 wire \heichips25_can_lehmann_fsm/net307 ;
 wire \heichips25_can_lehmann_fsm/net308 ;
 wire \heichips25_can_lehmann_fsm/net309 ;
 wire \heichips25_can_lehmann_fsm/net310 ;
 wire \heichips25_can_lehmann_fsm/net311 ;
 wire \heichips25_can_lehmann_fsm/net312 ;
 wire \heichips25_can_lehmann_fsm/net313 ;
 wire \heichips25_can_lehmann_fsm/net314 ;
 wire \heichips25_can_lehmann_fsm/net315 ;
 wire \heichips25_can_lehmann_fsm/net316 ;
 wire \heichips25_can_lehmann_fsm/net317 ;
 wire \heichips25_can_lehmann_fsm/net318 ;
 wire \heichips25_can_lehmann_fsm/net319 ;
 wire \heichips25_can_lehmann_fsm/net320 ;
 wire \heichips25_can_lehmann_fsm/net321 ;
 wire \heichips25_can_lehmann_fsm/net322 ;
 wire \heichips25_can_lehmann_fsm/net323 ;
 wire \heichips25_can_lehmann_fsm/net324 ;
 wire \heichips25_can_lehmann_fsm/net325 ;
 wire \heichips25_can_lehmann_fsm/net326 ;
 wire \heichips25_can_lehmann_fsm/net327 ;
 wire \heichips25_can_lehmann_fsm/net328 ;
 wire \heichips25_can_lehmann_fsm/net329 ;
 wire \heichips25_can_lehmann_fsm/net330 ;
 wire \heichips25_can_lehmann_fsm/net331 ;
 wire \heichips25_can_lehmann_fsm/net332 ;
 wire \heichips25_can_lehmann_fsm/net333 ;
 wire \heichips25_can_lehmann_fsm/net334 ;
 wire \heichips25_can_lehmann_fsm/net335 ;
 wire \heichips25_can_lehmann_fsm/net336 ;
 wire \heichips25_can_lehmann_fsm/net337 ;
 wire \heichips25_can_lehmann_fsm/net338 ;
 wire \heichips25_sap3/net339 ;
 wire \heichips25_sap3/net340 ;
 wire \heichips25_sap3/net341 ;
 wire \heichips25_sap3/net342 ;
 wire \heichips25_can_lehmann_fsm/net343 ;
 wire \heichips25_can_lehmann_fsm/net344 ;
 wire \heichips25_can_lehmann_fsm/net345 ;
 wire \heichips25_can_lehmann_fsm/net346 ;
 wire \heichips25_can_lehmann_fsm/net347 ;
 wire \heichips25_can_lehmann_fsm/net348 ;
 wire \heichips25_can_lehmann_fsm/net349 ;
 wire \heichips25_can_lehmann_fsm/net350 ;
 wire \heichips25_can_lehmann_fsm/net351 ;
 wire \heichips25_can_lehmann_fsm/net352 ;
 wire \heichips25_can_lehmann_fsm/net353 ;
 wire \heichips25_can_lehmann_fsm/net354 ;
 wire \heichips25_can_lehmann_fsm/net355 ;
 wire \heichips25_can_lehmann_fsm/net356 ;
 wire \heichips25_can_lehmann_fsm/net357 ;
 wire \heichips25_can_lehmann_fsm/net358 ;
 wire \heichips25_can_lehmann_fsm/net359 ;
 wire \heichips25_can_lehmann_fsm/net360 ;
 wire \heichips25_can_lehmann_fsm/net361 ;
 wire \heichips25_can_lehmann_fsm/net362 ;
 wire \heichips25_can_lehmann_fsm/net363 ;
 wire \heichips25_can_lehmann_fsm/net364 ;
 wire \heichips25_can_lehmann_fsm/net365 ;
 wire \heichips25_can_lehmann_fsm/net366 ;
 wire \heichips25_can_lehmann_fsm/net367 ;
 wire \heichips25_can_lehmann_fsm/net368 ;
 wire \heichips25_can_lehmann_fsm/net369 ;
 wire \heichips25_can_lehmann_fsm/net370 ;
 wire \heichips25_can_lehmann_fsm/net371 ;
 wire \heichips25_can_lehmann_fsm/net372 ;
 wire \heichips25_can_lehmann_fsm/net373 ;
 wire \heichips25_can_lehmann_fsm/net374 ;
 wire \heichips25_can_lehmann_fsm/net375 ;
 wire \heichips25_can_lehmann_fsm/net376 ;
 wire \heichips25_can_lehmann_fsm/net377 ;
 wire \heichips25_can_lehmann_fsm/net378 ;
 wire \heichips25_can_lehmann_fsm/net379 ;
 wire \heichips25_can_lehmann_fsm/net380 ;
 wire \heichips25_can_lehmann_fsm/net381 ;
 wire \heichips25_can_lehmann_fsm/net382 ;
 wire \heichips25_can_lehmann_fsm/net383 ;
 wire \heichips25_can_lehmann_fsm/net384 ;
 wire \heichips25_can_lehmann_fsm/net385 ;
 wire \heichips25_can_lehmann_fsm/net386 ;
 wire \heichips25_can_lehmann_fsm/net387 ;
 wire \heichips25_can_lehmann_fsm/net388 ;
 wire \heichips25_can_lehmann_fsm/net389 ;
 wire \heichips25_can_lehmann_fsm/net390 ;
 wire \heichips25_can_lehmann_fsm/net391 ;
 wire \heichips25_can_lehmann_fsm/net392 ;
 wire \heichips25_can_lehmann_fsm/net393 ;
 wire \heichips25_can_lehmann_fsm/net394 ;
 wire \heichips25_can_lehmann_fsm/net395 ;
 wire \heichips25_can_lehmann_fsm/net396 ;
 wire \heichips25_can_lehmann_fsm/net397 ;
 wire \heichips25_can_lehmann_fsm/net398 ;
 wire \heichips25_can_lehmann_fsm/net399 ;
 wire \heichips25_can_lehmann_fsm/net400 ;
 wire \heichips25_can_lehmann_fsm/net401 ;
 wire \heichips25_can_lehmann_fsm/net402 ;
 wire \heichips25_can_lehmann_fsm/net403 ;
 wire \heichips25_can_lehmann_fsm/net404 ;
 wire \heichips25_can_lehmann_fsm/net405 ;
 wire \heichips25_can_lehmann_fsm/net406 ;
 wire \heichips25_can_lehmann_fsm/net407 ;
 wire \heichips25_can_lehmann_fsm/net408 ;
 wire \heichips25_can_lehmann_fsm/net409 ;
 wire \heichips25_can_lehmann_fsm/net410 ;
 wire \heichips25_can_lehmann_fsm/net411 ;
 wire \heichips25_can_lehmann_fsm/net412 ;
 wire \heichips25_can_lehmann_fsm/net413 ;
 wire \heichips25_can_lehmann_fsm/net414 ;
 wire \heichips25_can_lehmann_fsm/net415 ;
 wire \heichips25_can_lehmann_fsm/net416 ;
 wire \heichips25_can_lehmann_fsm/net417 ;
 wire \heichips25_can_lehmann_fsm/net418 ;
 wire \heichips25_can_lehmann_fsm/net419 ;
 wire \heichips25_can_lehmann_fsm/net420 ;
 wire \heichips25_can_lehmann_fsm/net421 ;
 wire \heichips25_can_lehmann_fsm/net422 ;
 wire \heichips25_can_lehmann_fsm/net423 ;
 wire \heichips25_can_lehmann_fsm/net424 ;
 wire \heichips25_can_lehmann_fsm/net425 ;
 wire \heichips25_can_lehmann_fsm/net426 ;
 wire \heichips25_can_lehmann_fsm/net427 ;
 wire \heichips25_can_lehmann_fsm/net428 ;
 wire \heichips25_can_lehmann_fsm/net429 ;
 wire \heichips25_can_lehmann_fsm/net430 ;
 wire \heichips25_can_lehmann_fsm/net431 ;
 wire \heichips25_can_lehmann_fsm/net432 ;
 wire \heichips25_sap3/net433 ;
 wire \heichips25_sap3/net434 ;
 wire \heichips25_sap3/net435 ;
 wire \heichips25_sap3/net436 ;
 wire \heichips25_sap3/net437 ;
 wire \heichips25_sap3/net438 ;
 wire \heichips25_sap3/net439 ;
 wire \heichips25_sap3/net440 ;
 wire \heichips25_sap3/net441 ;
 wire \heichips25_sap3/net442 ;
 wire \heichips25_sap3/net443 ;
 wire \heichips25_sap3/net444 ;
 wire \heichips25_sap3/net445 ;
 wire \heichips25_sap3/net446 ;
 wire \heichips25_sap3/net447 ;
 wire \heichips25_sap3/net448 ;
 wire \heichips25_sap3/net449 ;
 wire \heichips25_sap3/net450 ;
 wire \heichips25_sap3/net451 ;
 wire \heichips25_sap3/net452 ;
 wire \heichips25_sap3/net453 ;
 wire \heichips25_sap3/net454 ;
 wire \heichips25_sap3/net455 ;
 wire \heichips25_sap3/net456 ;
 wire \heichips25_sap3/net457 ;
 wire \heichips25_sap3/net458 ;
 wire \heichips25_sap3/net459 ;
 wire \heichips25_sap3/net460 ;
 wire \heichips25_sap3/net461 ;
 wire \heichips25_sap3/net462 ;
 wire \heichips25_sap3/net463 ;
 wire \heichips25_can_lehmann_fsm/net464 ;
 wire \heichips25_can_lehmann_fsm/net465 ;
 wire \heichips25_can_lehmann_fsm/net466 ;
 wire \heichips25_can_lehmann_fsm/net467 ;
 wire \heichips25_can_lehmann_fsm/net468 ;
 wire \heichips25_can_lehmann_fsm/net469 ;
 wire \heichips25_can_lehmann_fsm/net470 ;
 wire \heichips25_can_lehmann_fsm/net471 ;
 wire \heichips25_can_lehmann_fsm/net472 ;
 wire \heichips25_can_lehmann_fsm/net473 ;
 wire \heichips25_can_lehmann_fsm/net474 ;
 wire \heichips25_can_lehmann_fsm/net475 ;
 wire \heichips25_can_lehmann_fsm/net476 ;
 wire \heichips25_can_lehmann_fsm/net477 ;
 wire \heichips25_can_lehmann_fsm/net478 ;
 wire \heichips25_can_lehmann_fsm/net479 ;
 wire \heichips25_can_lehmann_fsm/net480 ;
 wire \heichips25_can_lehmann_fsm/net481 ;
 wire \heichips25_can_lehmann_fsm/net482 ;
 wire \heichips25_can_lehmann_fsm/net483 ;
 wire \heichips25_can_lehmann_fsm/net484 ;
 wire \heichips25_can_lehmann_fsm/net485 ;
 wire \heichips25_can_lehmann_fsm/net486 ;
 wire \heichips25_can_lehmann_fsm/net487 ;
 wire \heichips25_can_lehmann_fsm/net488 ;
 wire \heichips25_can_lehmann_fsm/net489 ;
 wire \heichips25_can_lehmann_fsm/net490 ;
 wire \heichips25_can_lehmann_fsm/net491 ;
 wire \heichips25_can_lehmann_fsm/net492 ;
 wire \heichips25_can_lehmann_fsm/net493 ;
 wire \heichips25_can_lehmann_fsm/net494 ;
 wire \heichips25_can_lehmann_fsm/net495 ;
 wire \heichips25_can_lehmann_fsm/net496 ;
 wire \heichips25_can_lehmann_fsm/net497 ;
 wire \heichips25_can_lehmann_fsm/net498 ;
 wire \heichips25_can_lehmann_fsm/net499 ;
 wire \heichips25_can_lehmann_fsm/net500 ;
 wire \heichips25_can_lehmann_fsm/net501 ;
 wire \heichips25_can_lehmann_fsm/net502 ;
 wire \heichips25_can_lehmann_fsm/net503 ;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire \clknet_0_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_4_0_0_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_4_1_0_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_4_2_0_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_4_3_0_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_4_4_0_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_4_5_0_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_4_6_0_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_4_7_0_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_4_8_0_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_4_9_0_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_4_10_0_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_4_11_0_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_4_12_0_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_4_13_0_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_4_14_0_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_4_15_0_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_5_0__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_5_1__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_5_2__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_5_3__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_5_4__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_5_5__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_5_6__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_5_7__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_5_8__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_5_9__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_5_10__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_5_11__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_5_12__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_5_13__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_5_14__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_5_15__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_5_16__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_5_17__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_5_18__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_5_19__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_5_20__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_5_21__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_5_22__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_5_23__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_5_24__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_5_25__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_5_26__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_5_27__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_5_28__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_5_29__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_5_30__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \clknet_5_31__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ;
 wire \heichips25_sap3/net826 ;
 wire \heichips25_sap3/net827 ;
 wire \heichips25_sap3/net828 ;
 wire net829;
 wire \heichips25_sap3/net830 ;
 wire \heichips25_sap3/net831 ;
 wire \heichips25_sap3/net832 ;
 wire \heichips25_sap3/net833 ;
 wire \heichips25_sap3/clk_div_param_inst/net834 ;
 wire \heichips25_sap3/net835 ;
 wire \heichips25_sap3/net836 ;
 wire \heichips25_sap3/net837 ;
 wire \heichips25_sap3/net838 ;
 wire \heichips25_sap3/net839 ;
 wire \heichips25_can_lehmann_fsm/net840 ;
 wire \heichips25_can_lehmann_fsm/net841 ;
 wire \heichips25_can_lehmann_fsm/net842 ;
 wire \heichips25_can_lehmann_fsm/net843 ;
 wire \heichips25_can_lehmann_fsm/net844 ;
 wire \heichips25_can_lehmann_fsm/net845 ;
 wire \heichips25_can_lehmann_fsm/net846 ;
 wire \heichips25_can_lehmann_fsm/net847 ;
 wire \heichips25_can_lehmann_fsm/net848 ;
 wire \heichips25_can_lehmann_fsm/net849 ;
 wire \heichips25_can_lehmann_fsm/net850 ;
 wire \heichips25_can_lehmann_fsm/net851 ;
 wire \heichips25_can_lehmann_fsm/net852 ;
 wire \heichips25_can_lehmann_fsm/net853 ;
 wire \heichips25_can_lehmann_fsm/net854 ;
 wire \heichips25_can_lehmann_fsm/net855 ;
 wire \heichips25_can_lehmann_fsm/net856 ;
 wire \heichips25_can_lehmann_fsm/net857 ;
 wire \heichips25_can_lehmann_fsm/net858 ;
 wire \heichips25_can_lehmann_fsm/net859 ;
 wire \heichips25_can_lehmann_fsm/net860 ;
 wire \heichips25_can_lehmann_fsm/net861 ;
 wire \heichips25_can_lehmann_fsm/net862 ;
 wire \heichips25_can_lehmann_fsm/net863 ;
 wire \heichips25_can_lehmann_fsm/net864 ;
 wire \heichips25_can_lehmann_fsm/net865 ;
 wire \heichips25_can_lehmann_fsm/net866 ;
 wire \heichips25_can_lehmann_fsm/net867 ;
 wire \heichips25_can_lehmann_fsm/net868 ;
 wire \heichips25_can_lehmann_fsm/net869 ;
 wire \heichips25_can_lehmann_fsm/net870 ;
 wire \heichips25_can_lehmann_fsm/net871 ;
 wire \heichips25_can_lehmann_fsm/net872 ;
 wire \heichips25_can_lehmann_fsm/net873 ;
 wire \heichips25_can_lehmann_fsm/net874 ;
 wire \heichips25_can_lehmann_fsm/net875 ;
 wire \heichips25_can_lehmann_fsm/net876 ;
 wire \heichips25_can_lehmann_fsm/net877 ;
 wire \heichips25_can_lehmann_fsm/net878 ;
 wire \heichips25_can_lehmann_fsm/net879 ;
 wire \heichips25_can_lehmann_fsm/net880 ;
 wire \heichips25_can_lehmann_fsm/net881 ;
 wire \heichips25_can_lehmann_fsm/net882 ;
 wire \heichips25_can_lehmann_fsm/net883 ;
 wire \heichips25_can_lehmann_fsm/net884 ;
 wire \heichips25_can_lehmann_fsm/net885 ;
 wire \heichips25_can_lehmann_fsm/net886 ;
 wire \heichips25_can_lehmann_fsm/net887 ;
 wire \heichips25_can_lehmann_fsm/net888 ;
 wire \heichips25_can_lehmann_fsm/net889 ;
 wire \heichips25_can_lehmann_fsm/net890 ;
 wire \heichips25_sap3/net891 ;
 wire \heichips25_sap3/net892 ;
 wire \heichips25_can_lehmann_fsm/net893 ;
 wire \heichips25_can_lehmann_fsm/net894 ;
 wire \heichips25_can_lehmann_fsm/net895 ;
 wire \heichips25_can_lehmann_fsm/net896 ;
 wire \heichips25_can_lehmann_fsm/net897 ;
 wire \heichips25_can_lehmann_fsm/net898 ;
 wire \heichips25_can_lehmann_fsm/net899 ;
 wire \heichips25_can_lehmann_fsm/net900 ;
 wire \heichips25_can_lehmann_fsm/net901 ;
 wire \heichips25_can_lehmann_fsm/net902 ;
 wire \heichips25_can_lehmann_fsm/net903 ;
 wire \heichips25_can_lehmann_fsm/net904 ;
 wire \heichips25_can_lehmann_fsm/net905 ;
 wire \heichips25_can_lehmann_fsm/net906 ;
 wire \heichips25_can_lehmann_fsm/net907 ;
 wire \heichips25_can_lehmann_fsm/net908 ;
 wire \heichips25_can_lehmann_fsm/net909 ;
 wire \heichips25_can_lehmann_fsm/net910 ;
 wire \heichips25_can_lehmann_fsm/net911 ;
 wire \heichips25_can_lehmann_fsm/net912 ;
 wire \heichips25_can_lehmann_fsm/net913 ;
 wire \heichips25_can_lehmann_fsm/net914 ;
 wire \heichips25_can_lehmann_fsm/net915 ;
 wire \heichips25_can_lehmann_fsm/net916 ;
 wire \heichips25_can_lehmann_fsm/net917 ;
 wire \heichips25_can_lehmann_fsm/net918 ;
 wire \heichips25_can_lehmann_fsm/net919 ;
 wire \heichips25_can_lehmann_fsm/net920 ;
 wire \heichips25_can_lehmann_fsm/net921 ;
 wire \heichips25_can_lehmann_fsm/net922 ;
 wire \heichips25_can_lehmann_fsm/net923 ;
 wire \heichips25_can_lehmann_fsm/net924 ;
 wire \heichips25_sap3/net925 ;
 wire \heichips25_sap3/net926 ;
 wire \heichips25_can_lehmann_fsm/net927 ;
 wire \heichips25_can_lehmann_fsm/net928 ;
 wire \heichips25_can_lehmann_fsm/net929 ;
 wire \heichips25_can_lehmann_fsm/net930 ;
 wire \heichips25_can_lehmann_fsm/net931 ;
 wire \heichips25_can_lehmann_fsm/net932 ;
 wire \heichips25_can_lehmann_fsm/net933 ;
 wire \heichips25_can_lehmann_fsm/net934 ;
 wire \heichips25_can_lehmann_fsm/net935 ;
 wire \heichips25_can_lehmann_fsm/net936 ;
 wire \heichips25_can_lehmann_fsm/net937 ;
 wire \heichips25_can_lehmann_fsm/net938 ;
 wire \heichips25_can_lehmann_fsm/net939 ;
 wire \heichips25_can_lehmann_fsm/net940 ;
 wire \heichips25_can_lehmann_fsm/net941 ;
 wire \heichips25_can_lehmann_fsm/net942 ;
 wire \heichips25_can_lehmann_fsm/net943 ;
 wire \heichips25_can_lehmann_fsm/net944 ;
 wire \heichips25_can_lehmann_fsm/net945 ;
 wire \heichips25_can_lehmann_fsm/net946 ;
 wire \heichips25_can_lehmann_fsm/net947 ;
 wire \heichips25_can_lehmann_fsm/net948 ;
 wire \heichips25_can_lehmann_fsm/net949 ;
 wire \heichips25_can_lehmann_fsm/net950 ;
 wire \heichips25_can_lehmann_fsm/net951 ;
 wire \heichips25_can_lehmann_fsm/net952 ;
 wire \heichips25_sap3/net953 ;
 wire \heichips25_sap3/net954 ;
 wire \heichips25_can_lehmann_fsm/net955 ;
 wire \heichips25_can_lehmann_fsm/net956 ;
 wire \heichips25_can_lehmann_fsm/net957 ;
 wire \heichips25_can_lehmann_fsm/net958 ;
 wire \heichips25_can_lehmann_fsm/net959 ;
 wire \heichips25_can_lehmann_fsm/net960 ;
 wire \heichips25_can_lehmann_fsm/net961 ;
 wire \heichips25_can_lehmann_fsm/net962 ;
 wire \heichips25_can_lehmann_fsm/net963 ;
 wire \heichips25_can_lehmann_fsm/net964 ;
 wire \heichips25_can_lehmann_fsm/net965 ;
 wire \heichips25_can_lehmann_fsm/net966 ;
 wire \heichips25_can_lehmann_fsm/net967 ;
 wire \heichips25_can_lehmann_fsm/net968 ;
 wire \heichips25_can_lehmann_fsm/net969 ;
 wire \heichips25_can_lehmann_fsm/net970 ;
 wire \heichips25_can_lehmann_fsm/net971 ;
 wire \heichips25_can_lehmann_fsm/net972 ;
 wire \heichips25_can_lehmann_fsm/net973 ;
 wire \heichips25_can_lehmann_fsm/net974 ;
 wire \heichips25_can_lehmann_fsm/net975 ;
 wire \heichips25_can_lehmann_fsm/net976 ;
 wire \heichips25_can_lehmann_fsm/net977 ;
 wire \heichips25_can_lehmann_fsm/net978 ;
 wire \heichips25_can_lehmann_fsm/net979 ;
 wire \heichips25_can_lehmann_fsm/net980 ;
 wire \heichips25_can_lehmann_fsm/net981 ;
 wire \heichips25_can_lehmann_fsm/net982 ;
 wire \heichips25_can_lehmann_fsm/net983 ;
 wire \heichips25_can_lehmann_fsm/net984 ;
 wire \heichips25_can_lehmann_fsm/net985 ;
 wire \heichips25_can_lehmann_fsm/net986 ;
 wire \heichips25_can_lehmann_fsm/net987 ;
 wire \heichips25_can_lehmann_fsm/net988 ;
 wire \heichips25_can_lehmann_fsm/net989 ;
 wire \heichips25_can_lehmann_fsm/net990 ;
 wire \heichips25_can_lehmann_fsm/net991 ;
 wire \heichips25_can_lehmann_fsm/net992 ;
 wire \heichips25_can_lehmann_fsm/net993 ;
 wire \heichips25_can_lehmann_fsm/net994 ;
 wire \heichips25_can_lehmann_fsm/net995 ;
 wire \heichips25_can_lehmann_fsm/net996 ;
 wire \heichips25_can_lehmann_fsm/net997 ;
 wire \heichips25_can_lehmann_fsm/net998 ;
 wire \heichips25_can_lehmann_fsm/net999 ;
 wire \heichips25_can_lehmann_fsm/net1000 ;
 wire \heichips25_can_lehmann_fsm/net1001 ;
 wire \heichips25_can_lehmann_fsm/net1002 ;
 wire \heichips25_can_lehmann_fsm/net1003 ;
 wire \heichips25_can_lehmann_fsm/net1004 ;
 wire \heichips25_can_lehmann_fsm/net1005 ;
 wire \heichips25_can_lehmann_fsm/net1006 ;
 wire \heichips25_can_lehmann_fsm/net1007 ;
 wire \heichips25_can_lehmann_fsm/net1008 ;
 wire \heichips25_can_lehmann_fsm/net1009 ;
 wire \heichips25_can_lehmann_fsm/net1010 ;
 wire \heichips25_sap3/net1011 ;
 wire \heichips25_sap3/net1012 ;
 wire \heichips25_can_lehmann_fsm/net1013 ;
 wire \heichips25_can_lehmann_fsm/net1014 ;
 wire \heichips25_can_lehmann_fsm/net1015 ;
 wire \heichips25_can_lehmann_fsm/net1016 ;
 wire \heichips25_can_lehmann_fsm/net1017 ;
 wire \heichips25_can_lehmann_fsm/net1018 ;
 wire \heichips25_sap3/net1019 ;
 wire \heichips25_sap3/net1020 ;
 wire \heichips25_can_lehmann_fsm/net1021 ;
 wire \heichips25_can_lehmann_fsm/net1022 ;
 wire \heichips25_can_lehmann_fsm/net1023 ;
 wire \heichips25_can_lehmann_fsm/net1024 ;
 wire \heichips25_can_lehmann_fsm/net1025 ;
 wire \heichips25_can_lehmann_fsm/net1026 ;
 wire \heichips25_can_lehmann_fsm/net1027 ;
 wire \heichips25_can_lehmann_fsm/net1028 ;
 wire \heichips25_can_lehmann_fsm/net1029 ;
 wire \heichips25_can_lehmann_fsm/net1030 ;
 wire \heichips25_sap3/net1031 ;
 wire \heichips25_sap3/net1032 ;
 wire \heichips25_can_lehmann_fsm/net1033 ;
 wire \heichips25_can_lehmann_fsm/net1034 ;
 wire \heichips25_can_lehmann_fsm/net1035 ;
 wire \heichips25_can_lehmann_fsm/net1036 ;
 wire \heichips25_can_lehmann_fsm/net1037 ;
 wire \heichips25_can_lehmann_fsm/net1038 ;
 wire \heichips25_can_lehmann_fsm/net1039 ;
 wire \heichips25_can_lehmann_fsm/net1040 ;
 wire \heichips25_can_lehmann_fsm/net1041 ;
 wire \heichips25_can_lehmann_fsm/net1042 ;
 wire \heichips25_can_lehmann_fsm/net1043 ;
 wire \heichips25_can_lehmann_fsm/net1044 ;
 wire \heichips25_can_lehmann_fsm/net1045 ;
 wire \heichips25_can_lehmann_fsm/net1046 ;
 wire \heichips25_can_lehmann_fsm/net1047 ;
 wire \heichips25_can_lehmann_fsm/net1048 ;
 wire \heichips25_can_lehmann_fsm/net1049 ;
 wire \heichips25_can_lehmann_fsm/net1050 ;
 wire \heichips25_can_lehmann_fsm/net1051 ;
 wire \heichips25_can_lehmann_fsm/net1052 ;
 wire \heichips25_can_lehmann_fsm/net1053 ;
 wire \heichips25_can_lehmann_fsm/net1054 ;
 wire \heichips25_can_lehmann_fsm/net1055 ;
 wire \heichips25_can_lehmann_fsm/net1056 ;
 wire \heichips25_can_lehmann_fsm/net1057 ;
 wire \heichips25_sap3/net1058 ;
 wire \heichips25_sap3/net1059 ;
 wire \heichips25_can_lehmann_fsm/net1060 ;
 wire \heichips25_can_lehmann_fsm/net1061 ;
 wire \heichips25_can_lehmann_fsm/net1062 ;
 wire \heichips25_can_lehmann_fsm/net1063 ;
 wire \heichips25_sap3/net1064 ;
 wire \heichips25_sap3/net1065 ;
 wire \heichips25_can_lehmann_fsm/net1066 ;
 wire \heichips25_can_lehmann_fsm/net1067 ;
 wire \heichips25_can_lehmann_fsm/net1068 ;
 wire \heichips25_can_lehmann_fsm/net1069 ;
 wire \heichips25_can_lehmann_fsm/net1070 ;
 wire \heichips25_sap3/net1071 ;
 wire \heichips25_sap3/net1072 ;
 wire \heichips25_sap3/net1073 ;
 wire \heichips25_can_lehmann_fsm/net1074 ;
 wire \heichips25_can_lehmann_fsm/net1075 ;
 wire \heichips25_can_lehmann_fsm/net1076 ;
 wire \heichips25_can_lehmann_fsm/net1077 ;
 wire \heichips25_can_lehmann_fsm/net1078 ;
 wire \heichips25_can_lehmann_fsm/net1079 ;
 wire \heichips25_can_lehmann_fsm/net1080 ;
 wire \heichips25_can_lehmann_fsm/net1081 ;
 wire \heichips25_can_lehmann_fsm/net1082 ;
 wire \heichips25_can_lehmann_fsm/net1083 ;
 wire \heichips25_can_lehmann_fsm/net1084 ;
 wire \heichips25_can_lehmann_fsm/net1085 ;
 wire \heichips25_can_lehmann_fsm/net1086 ;
 wire \heichips25_can_lehmann_fsm/net1087 ;
 wire \heichips25_can_lehmann_fsm/net1088 ;
 wire \heichips25_can_lehmann_fsm/net1089 ;
 wire \heichips25_can_lehmann_fsm/net1090 ;
 wire \heichips25_can_lehmann_fsm/net1091 ;
 wire \heichips25_can_lehmann_fsm/net1092 ;
 wire \heichips25_can_lehmann_fsm/net1093 ;
 wire \heichips25_can_lehmann_fsm/net1094 ;
 wire \heichips25_can_lehmann_fsm/net1095 ;
 wire \heichips25_can_lehmann_fsm/net1096 ;
 wire \heichips25_can_lehmann_fsm/net1097 ;
 wire \heichips25_can_lehmann_fsm/net1098 ;
 wire \heichips25_can_lehmann_fsm/net1099 ;
 wire \heichips25_can_lehmann_fsm/net1100 ;
 wire \heichips25_can_lehmann_fsm/net1101 ;
 wire \heichips25_can_lehmann_fsm/net1102 ;
 wire \heichips25_can_lehmann_fsm/net1103 ;
 wire \heichips25_can_lehmann_fsm/net1104 ;
 wire \heichips25_sap3/net1105 ;
 wire \heichips25_can_lehmann_fsm/net1106 ;
 wire \heichips25_can_lehmann_fsm/net1107 ;
 wire \heichips25_can_lehmann_fsm/net1108 ;
 wire \heichips25_can_lehmann_fsm/net1109 ;
 wire \heichips25_can_lehmann_fsm/net1110 ;
 wire \heichips25_can_lehmann_fsm/net1111 ;
 wire \heichips25_sap3/net1112 ;
 wire \heichips25_can_lehmann_fsm/net1113 ;
 wire \heichips25_can_lehmann_fsm/net1114 ;
 wire \heichips25_can_lehmann_fsm/net1115 ;
 wire \heichips25_can_lehmann_fsm/net1116 ;
 wire \heichips25_can_lehmann_fsm/net1117 ;
 wire \heichips25_can_lehmann_fsm/net1118 ;
 wire \heichips25_sap3/net1119 ;
 wire \heichips25_sap3/net1120 ;
 wire \heichips25_sap3/net1121 ;
 wire \heichips25_can_lehmann_fsm/net1122 ;
 wire \heichips25_can_lehmann_fsm/net1123 ;
 wire \heichips25_sap3/net1124 ;
 wire \heichips25_sap3/net1125 ;
 wire \heichips25_can_lehmann_fsm/net1126 ;
 wire \heichips25_can_lehmann_fsm/net1127 ;
 wire \heichips25_sap3/net1128 ;
 wire \heichips25_can_lehmann_fsm/net1129 ;
 wire \heichips25_sap3/net1130 ;
 wire \heichips25_sap3/net1131 ;
 wire \heichips25_can_lehmann_fsm/net1132 ;
 wire \heichips25_can_lehmann_fsm/net1133 ;
 wire \heichips25_can_lehmann_fsm/net1134 ;
 wire \heichips25_can_lehmann_fsm/net1135 ;
 wire \heichips25_can_lehmann_fsm/net1136 ;
 wire \heichips25_can_lehmann_fsm/net1137 ;
 wire \heichips25_sap3/net1138 ;
 wire \heichips25_can_lehmann_fsm/net1139 ;
 wire \heichips25_can_lehmann_fsm/net1140 ;
 wire \heichips25_sap3/net1141 ;
 wire \heichips25_can_lehmann_fsm/net1142 ;
 wire \heichips25_sap3/net1143 ;
 wire \heichips25_sap3/net1144 ;
 wire \heichips25_sap3/net1145 ;
 wire \heichips25_can_lehmann_fsm/net1146 ;
 wire \heichips25_can_lehmann_fsm/net1147 ;
 wire \heichips25_can_lehmann_fsm/net1148 ;
 wire \heichips25_sap3/net1149 ;
 wire \heichips25_can_lehmann_fsm/net1150 ;
 wire \heichips25_can_lehmann_fsm/net1151 ;
 wire \heichips25_can_lehmann_fsm/net1152 ;
 wire \heichips25_can_lehmann_fsm/net1153 ;
 wire \heichips25_can_lehmann_fsm/net1154 ;
 wire \heichips25_can_lehmann_fsm/net1155 ;
 wire \heichips25_can_lehmann_fsm/net1156 ;
 wire \heichips25_can_lehmann_fsm/net1157 ;
 wire \heichips25_can_lehmann_fsm/net1158 ;
 wire \heichips25_can_lehmann_fsm/net1159 ;
 wire \heichips25_can_lehmann_fsm/net1160 ;
 wire \heichips25_can_lehmann_fsm/net1161 ;
 wire \heichips25_sap3/net1162 ;
 wire \heichips25_sap3/net1163 ;
 wire \heichips25_can_lehmann_fsm/net1164 ;
 wire \heichips25_can_lehmann_fsm/net1165 ;
 wire \heichips25_can_lehmann_fsm/net1166 ;
 wire \heichips25_can_lehmann_fsm/net1167 ;
 wire \heichips25_can_lehmann_fsm/net1168 ;
 wire \heichips25_can_lehmann_fsm/net1169 ;
 wire \heichips25_can_lehmann_fsm/net1170 ;
 wire \heichips25_can_lehmann_fsm/net1171 ;
 wire \heichips25_can_lehmann_fsm/net1172 ;
 wire \heichips25_can_lehmann_fsm/net1173 ;
 wire \heichips25_can_lehmann_fsm/net1174 ;
 wire \heichips25_can_lehmann_fsm/net1175 ;
 wire \heichips25_sap3/net1176 ;
 wire \heichips25_can_lehmann_fsm/net1177 ;
 wire \heichips25_sap3/net1178 ;
 wire \heichips25_sap3/net1179 ;
 wire \heichips25_can_lehmann_fsm/net1180 ;
 wire \heichips25_can_lehmann_fsm/net1181 ;
 wire \heichips25_can_lehmann_fsm/net1182 ;
 wire \heichips25_can_lehmann_fsm/net1183 ;
 wire \heichips25_can_lehmann_fsm/net1184 ;
 wire \heichips25_can_lehmann_fsm/net1185 ;
 wire \heichips25_can_lehmann_fsm/net1186 ;
 wire \heichips25_can_lehmann_fsm/net1187 ;
 wire \heichips25_can_lehmann_fsm/net1188 ;
 wire \heichips25_can_lehmann_fsm/net1189 ;
 wire \heichips25_can_lehmann_fsm/net1190 ;
 wire \heichips25_can_lehmann_fsm/net1191 ;
 wire \heichips25_can_lehmann_fsm/net1192 ;
 wire \heichips25_can_lehmann_fsm/net1193 ;
 wire \heichips25_can_lehmann_fsm/net1194 ;
 wire \heichips25_can_lehmann_fsm/net1195 ;
 wire \heichips25_can_lehmann_fsm/net1196 ;
 wire \heichips25_sap3/net1197 ;
 wire \heichips25_can_lehmann_fsm/net1198 ;
 wire \heichips25_can_lehmann_fsm/net1199 ;
 wire \heichips25_can_lehmann_fsm/net1200 ;
 wire \heichips25_can_lehmann_fsm/net1201 ;
 wire \heichips25_can_lehmann_fsm/net1202 ;
 wire \heichips25_can_lehmann_fsm/net1203 ;
 wire \heichips25_can_lehmann_fsm/net1204 ;
 wire \heichips25_can_lehmann_fsm/net1205 ;
 wire \heichips25_can_lehmann_fsm/net1206 ;
 wire \heichips25_can_lehmann_fsm/net1207 ;
 wire \heichips25_can_lehmann_fsm/net1208 ;
 wire \heichips25_can_lehmann_fsm/net1209 ;
 wire \heichips25_can_lehmann_fsm/net1210 ;
 wire \heichips25_can_lehmann_fsm/net1211 ;
 wire \heichips25_can_lehmann_fsm/net1212 ;
 wire \heichips25_can_lehmann_fsm/net1213 ;
 wire \heichips25_can_lehmann_fsm/net1214 ;
 wire \heichips25_can_lehmann_fsm/net1215 ;
 wire \heichips25_can_lehmann_fsm/net1216 ;
 wire \heichips25_can_lehmann_fsm/net1217 ;
 wire \heichips25_can_lehmann_fsm/net1218 ;
 wire \heichips25_can_lehmann_fsm/net1219 ;
 wire \heichips25_can_lehmann_fsm/net1220 ;
 wire \heichips25_can_lehmann_fsm/net1221 ;
 wire \heichips25_can_lehmann_fsm/net1222 ;
 wire \heichips25_sap3/net1223 ;
 wire \heichips25_sap3/net1224 ;
 wire \heichips25_sap3/net1225 ;
 wire \heichips25_can_lehmann_fsm/net1226 ;
 wire \heichips25_can_lehmann_fsm/net1227 ;
 wire \heichips25_can_lehmann_fsm/net1228 ;
 wire \heichips25_can_lehmann_fsm/net1229 ;
 wire \heichips25_can_lehmann_fsm/net1230 ;
 wire \heichips25_can_lehmann_fsm/net1231 ;
 wire \heichips25_can_lehmann_fsm/net1232 ;
 wire \heichips25_can_lehmann_fsm/net1233 ;
 wire \heichips25_can_lehmann_fsm/net1234 ;
 wire \heichips25_can_lehmann_fsm/net1235 ;
 wire \heichips25_can_lehmann_fsm/net1236 ;
 wire \heichips25_can_lehmann_fsm/net1237 ;
 wire \heichips25_can_lehmann_fsm/net1238 ;
 wire \heichips25_can_lehmann_fsm/net1239 ;
 wire \heichips25_can_lehmann_fsm/net1240 ;
 wire \heichips25_can_lehmann_fsm/net1241 ;
 wire \heichips25_can_lehmann_fsm/net1242 ;
 wire \heichips25_can_lehmann_fsm/net1243 ;
 wire \heichips25_can_lehmann_fsm/net1244 ;
 wire \heichips25_can_lehmann_fsm/net1245 ;
 wire \heichips25_can_lehmann_fsm/net1246 ;
 wire \heichips25_can_lehmann_fsm/net1247 ;
 wire \heichips25_can_lehmann_fsm/net1248 ;
 wire \heichips25_can_lehmann_fsm/net1249 ;
 wire \heichips25_can_lehmann_fsm/net1250 ;
 wire \heichips25_can_lehmann_fsm/net1251 ;
 wire \heichips25_can_lehmann_fsm/net1252 ;
 wire \heichips25_can_lehmann_fsm/net1253 ;
 wire \heichips25_can_lehmann_fsm/net1254 ;
 wire \heichips25_can_lehmann_fsm/net1255 ;
 wire \heichips25_can_lehmann_fsm/net1256 ;
 wire \heichips25_can_lehmann_fsm/net1257 ;
 wire \heichips25_can_lehmann_fsm/net1258 ;
 wire \heichips25_can_lehmann_fsm/net1259 ;
 wire \heichips25_can_lehmann_fsm/net1260 ;
 wire \heichips25_can_lehmann_fsm/net1261 ;
 wire \heichips25_can_lehmann_fsm/net1262 ;
 wire \heichips25_can_lehmann_fsm/net1263 ;
 wire \heichips25_can_lehmann_fsm/net1264 ;
 wire \heichips25_can_lehmann_fsm/net1265 ;
 wire \heichips25_can_lehmann_fsm/net1266 ;
 wire \heichips25_can_lehmann_fsm/net1267 ;
 wire \heichips25_can_lehmann_fsm/net1268 ;
 wire \heichips25_can_lehmann_fsm/net1269 ;
 wire \heichips25_can_lehmann_fsm/net1270 ;
 wire \heichips25_can_lehmann_fsm/net1271 ;
 wire \heichips25_can_lehmann_fsm/net1272 ;
 wire \heichips25_can_lehmann_fsm/net1273 ;
 wire \heichips25_can_lehmann_fsm/net1274 ;
 wire \heichips25_sap3/net1275 ;
 wire \heichips25_sap3/net1276 ;
 wire \heichips25_can_lehmann_fsm/net1277 ;
 wire \heichips25_can_lehmann_fsm/net1278 ;
 wire \heichips25_can_lehmann_fsm/net1279 ;

 sg13g2_nor2b_1 _04_ (.A(net507),
    .B_N(net2),
    .Y(_00_));
 sg13g2_and2_1 _05_ (.A(net2),
    .B(net1),
    .X(_01_));
 sg13g2_mux2_1 _06_ (.A0(\uo_out_fsm[0] ),
    .A1(\uo_out_sap3[0] ),
    .S(net507),
    .X(net35));
 sg13g2_mux2_1 _07_ (.A0(\uo_out_fsm[1] ),
    .A1(\uo_out_sap3[1] ),
    .S(net504),
    .X(net36));
 sg13g2_mux2_1 _08_ (.A0(\uo_out_fsm[2] ),
    .A1(\uo_out_sap3[2] ),
    .S(net507),
    .X(net37));
 sg13g2_mux2_1 _09_ (.A0(\uo_out_fsm[3] ),
    .A1(\uo_out_sap3[3] ),
    .S(net507),
    .X(net38));
 sg13g2_mux2_1 _10_ (.A0(\uo_out_fsm[4] ),
    .A1(\uo_out_sap3[4] ),
    .S(net507),
    .X(net39));
 sg13g2_mux2_1 _11_ (.A0(\uo_out_fsm[5] ),
    .A1(\uo_out_sap3[5] ),
    .S(net507),
    .X(net40));
 sg13g2_mux2_1 _12_ (.A0(\uo_out_fsm[6] ),
    .A1(net523),
    .S(net507),
    .X(net41));
 sg13g2_mux2_1 _13_ (.A0(\uo_out_fsm[7] ),
    .A1(net524),
    .S(net507),
    .X(net42));
 sg13g2_mux2_1 _14_ (.A0(net515),
    .A1(\uio_out_sap3[0] ),
    .S(net504),
    .X(net27));
 sg13g2_mux2_1 _15_ (.A0(net516),
    .A1(\uio_out_sap3[1] ),
    .S(net504),
    .X(net28));
 sg13g2_mux2_1 _16_ (.A0(net517),
    .A1(net44),
    .S(net504),
    .X(net29));
 sg13g2_mux2_1 _17_ (.A0(net518),
    .A1(\uio_out_sap3[3] ),
    .S(net504),
    .X(net30));
 sg13g2_mux2_1 _18_ (.A0(net519),
    .A1(net46),
    .S(net504),
    .X(net31));
 sg13g2_mux2_1 _19_ (.A0(net520),
    .A1(\uio_out_sap3[5] ),
    .S(net504),
    .X(net32));
 sg13g2_mux2_1 _20_ (.A0(net521),
    .A1(net43),
    .S(net504),
    .X(net33));
 sg13g2_mux2_1 _21_ (.A0(net522),
    .A1(net47),
    .S(net505),
    .X(net34));
 sg13g2_mux2_1 _22_ (.A0(net),
    .A1(\uio_oe_sap3[0] ),
    .S(net505),
    .X(net19));
 sg13g2_mux2_1 _23_ (.A0(net508),
    .A1(\uio_oe_sap3[1] ),
    .S(net505),
    .X(net20));
 sg13g2_mux2_1 _24_ (.A0(net509),
    .A1(\uio_oe_sap3[2] ),
    .S(net505),
    .X(net21));
 sg13g2_mux2_1 _25_ (.A0(net510),
    .A1(\uio_oe_sap3[3] ),
    .S(net506),
    .X(net22));
 sg13g2_mux2_1 _26_ (.A0(net511),
    .A1(\uio_oe_sap3[4] ),
    .S(net506),
    .X(net23));
 sg13g2_mux2_1 _27_ (.A0(net512),
    .A1(net829),
    .S(net506),
    .X(net24));
 sg13g2_mux2_1 _28_ (.A0(net513),
    .A1(\uio_oe_sap3[6] ),
    .S(net506),
    .X(net25));
 sg13g2_mux2_1 _29_ (.A0(net514),
    .A1(\uio_oe_sap3[7] ),
    .S(net506),
    .X(net26));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3061__526  (.L_HI(net525));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1528_  (.Y(\heichips25_can_lehmann_fsm/_0852_ ),
    .A(\heichips25_can_lehmann_fsm/net1132 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1529_  (.Y(\heichips25_can_lehmann_fsm/_0853_ ),
    .A(\heichips25_can_lehmann_fsm/net1142 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1530_  (.Y(\heichips25_can_lehmann_fsm/_0854_ ),
    .A(\heichips25_can_lehmann_fsm/net1043 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1531_  (.Y(\heichips25_can_lehmann_fsm/_0855_ ),
    .A(\heichips25_can_lehmann_fsm/net1051 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1532_  (.Y(\heichips25_can_lehmann_fsm/_0856_ ),
    .A(\heichips25_can_lehmann_fsm/net1155 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1533_  (.Y(\heichips25_can_lehmann_fsm/_0857_ ),
    .A(\heichips25_can_lehmann_fsm/net1117 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1534_  (.Y(\heichips25_can_lehmann_fsm/_0858_ ),
    .A(\heichips25_can_lehmann_fsm/net1147 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1535_  (.Y(\heichips25_can_lehmann_fsm/_0859_ ),
    .A(\heichips25_can_lehmann_fsm/net1151 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1536_  (.Y(\heichips25_can_lehmann_fsm/_0860_ ),
    .A(\heichips25_can_lehmann_fsm/net1229 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1537_  (.Y(\heichips25_can_lehmann_fsm/_0861_ ),
    .A(\heichips25_can_lehmann_fsm/net877 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1538_  (.Y(\heichips25_can_lehmann_fsm/_0862_ ),
    .A(\heichips25_can_lehmann_fsm/net944 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1539_  (.Y(\heichips25_can_lehmann_fsm/_0863_ ),
    .A(\heichips25_can_lehmann_fsm/net842 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1540_  (.Y(\heichips25_can_lehmann_fsm/_0864_ ),
    .A(\heichips25_can_lehmann_fsm/net1164 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1541_  (.Y(\heichips25_can_lehmann_fsm/_0865_ ),
    .A(\heichips25_can_lehmann_fsm/net1160 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1542_  (.Y(\heichips25_can_lehmann_fsm/_0866_ ),
    .A(\heichips25_can_lehmann_fsm/net993 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1543_  (.Y(\heichips25_can_lehmann_fsm/_0867_ ),
    .A(\heichips25_can_lehmann_fsm/net951 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1544_  (.Y(\heichips25_can_lehmann_fsm/_0868_ ),
    .A(\heichips25_can_lehmann_fsm/net1152 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1545_  (.Y(\heichips25_can_lehmann_fsm/_0869_ ),
    .A(\heichips25_can_lehmann_fsm/net960 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1546_  (.Y(\heichips25_can_lehmann_fsm/_0870_ ),
    .A(\heichips25_can_lehmann_fsm/net1074 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1547_  (.Y(\heichips25_can_lehmann_fsm/_0871_ ),
    .A(\heichips25_can_lehmann_fsm/net849 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1548_  (.Y(\heichips25_can_lehmann_fsm/_0872_ ),
    .A(\heichips25_can_lehmann_fsm/net1146 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1549_  (.Y(\heichips25_can_lehmann_fsm/_0873_ ),
    .A(\heichips25_can_lehmann_fsm/net990 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1550_  (.Y(\heichips25_can_lehmann_fsm/_0874_ ),
    .A(\heichips25_can_lehmann_fsm/net998 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1551_  (.Y(\heichips25_can_lehmann_fsm/_0875_ ),
    .A(\heichips25_can_lehmann_fsm/net853 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1552_  (.Y(\heichips25_can_lehmann_fsm/_0876_ ),
    .A(\heichips25_can_lehmann_fsm/net1129 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1553_  (.Y(\heichips25_can_lehmann_fsm/_0877_ ),
    .A(\heichips25_can_lehmann_fsm/net881 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1554_  (.Y(\heichips25_can_lehmann_fsm/_0878_ ),
    .A(\heichips25_can_lehmann_fsm/net867 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1555_  (.Y(\heichips25_can_lehmann_fsm/_0879_ ),
    .A(\heichips25_can_lehmann_fsm/net1139 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1556_  (.Y(\heichips25_can_lehmann_fsm/_0880_ ),
    .A(\heichips25_can_lehmann_fsm/net931 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1557_  (.Y(\heichips25_can_lehmann_fsm/_0881_ ),
    .A(\heichips25_can_lehmann_fsm/net906 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1558_  (.Y(\heichips25_can_lehmann_fsm/_0882_ ),
    .A(\heichips25_can_lehmann_fsm/net1122 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1559_  (.Y(\heichips25_can_lehmann_fsm/_0883_ ),
    .A(\heichips25_can_lehmann_fsm/net844 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1560_  (.Y(\heichips25_can_lehmann_fsm/_0884_ ),
    .A(\heichips25_can_lehmann_fsm/net860 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1561_  (.Y(\heichips25_can_lehmann_fsm/_0885_ ),
    .A(\heichips25_can_lehmann_fsm/net855 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1562_  (.Y(\heichips25_can_lehmann_fsm/_0886_ ),
    .A(\heichips25_can_lehmann_fsm/net1090 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1563_  (.Y(\heichips25_can_lehmann_fsm/_0887_ ),
    .A(\heichips25_can_lehmann_fsm/net928 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1564_  (.Y(\heichips25_can_lehmann_fsm/_0888_ ),
    .A(\heichips25_can_lehmann_fsm/net995 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1565_  (.Y(\heichips25_can_lehmann_fsm/_0889_ ),
    .A(\heichips25_can_lehmann_fsm/net918 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1566_  (.Y(\heichips25_can_lehmann_fsm/_0890_ ),
    .A(\heichips25_can_lehmann_fsm/net1021 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1567_  (.Y(\heichips25_can_lehmann_fsm/_0891_ ),
    .A(\heichips25_can_lehmann_fsm/net889 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1568_  (.Y(\heichips25_can_lehmann_fsm/_0892_ ),
    .A(\heichips25_can_lehmann_fsm/net978 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1569_  (.Y(\heichips25_can_lehmann_fsm/_0893_ ),
    .A(\heichips25_can_lehmann_fsm/net985 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1570_  (.Y(\heichips25_can_lehmann_fsm/_0894_ ),
    .A(\heichips25_can_lehmann_fsm/net1022 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1571_  (.Y(\heichips25_can_lehmann_fsm/_0895_ ),
    .A(\heichips25_can_lehmann_fsm/net872 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1572_  (.Y(\heichips25_can_lehmann_fsm/_0896_ ),
    .A(\heichips25_can_lehmann_fsm/net927 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1573_  (.Y(\heichips25_can_lehmann_fsm/_0897_ ),
    .A(\heichips25_can_lehmann_fsm/net846 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1574_  (.Y(\heichips25_can_lehmann_fsm/_0898_ ),
    .A(\heichips25_can_lehmann_fsm/net957 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1575_  (.Y(\heichips25_can_lehmann_fsm/_0899_ ),
    .A(\heichips25_can_lehmann_fsm/net946 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1576_  (.Y(\heichips25_can_lehmann_fsm/_0900_ ),
    .A(\heichips25_can_lehmann_fsm/net887 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1577_  (.Y(\heichips25_can_lehmann_fsm/_0901_ ),
    .A(\heichips25_can_lehmann_fsm/net885 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1578_  (.Y(\heichips25_can_lehmann_fsm/_0902_ ),
    .A(\heichips25_can_lehmann_fsm/net874 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1579_  (.Y(\heichips25_can_lehmann_fsm/_0903_ ),
    .A(\heichips25_can_lehmann_fsm/net1083 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1580_  (.Y(\heichips25_can_lehmann_fsm/_0904_ ),
    .A(\heichips25_can_lehmann_fsm/net1017 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1581_  (.Y(\heichips25_can_lehmann_fsm/_0905_ ),
    .A(\heichips25_can_lehmann_fsm/net1045 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1582_  (.Y(\heichips25_can_lehmann_fsm/_0906_ ),
    .A(\heichips25_can_lehmann_fsm/net1035 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1583_  (.Y(\heichips25_can_lehmann_fsm/_0907_ ),
    .A(\heichips25_can_lehmann_fsm/net1027 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1584_  (.Y(\heichips25_can_lehmann_fsm/_0908_ ),
    .A(\heichips25_can_lehmann_fsm/net1103 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1585_  (.Y(\heichips25_can_lehmann_fsm/_0909_ ),
    .A(\heichips25_can_lehmann_fsm/net1077 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1586_  (.Y(\heichips25_can_lehmann_fsm/_0910_ ),
    .A(\heichips25_can_lehmann_fsm/net1060 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1587_  (.Y(\heichips25_can_lehmann_fsm/_0911_ ),
    .A(\heichips25_can_lehmann_fsm/net934 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1588_  (.Y(\heichips25_can_lehmann_fsm/_0912_ ),
    .A(\heichips25_can_lehmann_fsm/net904 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1589_  (.Y(\heichips25_can_lehmann_fsm/_0913_ ),
    .A(\heichips25_can_lehmann_fsm/net1025 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1590_  (.Y(\heichips25_can_lehmann_fsm/_0914_ ),
    .A(\heichips25_can_lehmann_fsm/net970 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1591_  (.Y(\heichips25_can_lehmann_fsm/_0915_ ),
    .A(\heichips25_can_lehmann_fsm/net1097 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1592_  (.Y(\heichips25_can_lehmann_fsm/_0916_ ),
    .A(\heichips25_can_lehmann_fsm/net1013 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1593_  (.Y(\heichips25_can_lehmann_fsm/_0917_ ),
    .A(\heichips25_can_lehmann_fsm/net1106 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1594_  (.Y(\heichips25_can_lehmann_fsm/_0918_ ),
    .A(\heichips25_can_lehmann_fsm/net863 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1595_  (.Y(\heichips25_can_lehmann_fsm/_0919_ ),
    .A(\heichips25_can_lehmann_fsm/net992 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1596_  (.Y(\heichips25_can_lehmann_fsm/_0920_ ),
    .A(\heichips25_can_lehmann_fsm/net858 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1597_  (.Y(\heichips25_can_lehmann_fsm/_0921_ ),
    .A(\heichips25_can_lehmann_fsm/net1062 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1598_  (.Y(\heichips25_can_lehmann_fsm/_0922_ ),
    .A(\heichips25_can_lehmann_fsm/net1047 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1599_  (.Y(\heichips25_can_lehmann_fsm/_0923_ ),
    .A(\heichips25_can_lehmann_fsm/net893 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1600_  (.Y(\heichips25_can_lehmann_fsm/_0924_ ),
    .A(\heichips25_can_lehmann_fsm/net937 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1601_  (.Y(\heichips25_can_lehmann_fsm/_0925_ ),
    .A(\heichips25_can_lehmann_fsm/net981 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1602_  (.Y(\heichips25_can_lehmann_fsm/_0926_ ),
    .A(\heichips25_can_lehmann_fsm/net1108 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1603_  (.Y(\heichips25_can_lehmann_fsm/_0927_ ),
    .A(\heichips25_can_lehmann_fsm/net861 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1604_  (.Y(\heichips25_can_lehmann_fsm/_0928_ ),
    .A(\heichips25_can_lehmann_fsm/net1049 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1605_  (.Y(\heichips25_can_lehmann_fsm/_0929_ ),
    .A(\heichips25_can_lehmann_fsm/net966 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1606_  (.Y(\heichips25_can_lehmann_fsm/_0930_ ),
    .A(\heichips25_can_lehmann_fsm/net909 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1607_  (.Y(\heichips25_can_lehmann_fsm/_0931_ ),
    .A(\heichips25_can_lehmann_fsm/net900 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1608_  (.Y(\heichips25_can_lehmann_fsm/_0932_ ),
    .A(\heichips25_can_lehmann_fsm/net1041 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1609_  (.Y(\heichips25_can_lehmann_fsm/_0933_ ),
    .A(\heichips25_can_lehmann_fsm/net996 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1610_  (.Y(\heichips25_can_lehmann_fsm/_0934_ ),
    .A(\heichips25_can_lehmann_fsm/net1008 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1611_  (.Y(\heichips25_can_lehmann_fsm/_0935_ ),
    .A(\heichips25_can_lehmann_fsm/net1056 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1612_  (.Y(\heichips25_can_lehmann_fsm/_0936_ ),
    .A(\heichips25_can_lehmann_fsm/net913 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1613_  (.Y(\heichips25_can_lehmann_fsm/_0937_ ),
    .A(\heichips25_can_lehmann_fsm/net865 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1614_  (.Y(\heichips25_can_lehmann_fsm/_0938_ ),
    .A(\heichips25_can_lehmann_fsm/net1100 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1615_  (.Y(\heichips25_can_lehmann_fsm/_0939_ ),
    .A(\heichips25_can_lehmann_fsm/net955 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1616_  (.Y(\heichips25_can_lehmann_fsm/_0940_ ),
    .A(\heichips25_can_lehmann_fsm/net870 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1617_  (.Y(\heichips25_can_lehmann_fsm/_0941_ ),
    .A(\heichips25_can_lehmann_fsm/net1003 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1618_  (.Y(\heichips25_can_lehmann_fsm/_0942_ ),
    .A(\heichips25_can_lehmann_fsm/net1177 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1619_  (.Y(\heichips25_can_lehmann_fsm/_0943_ ),
    .A(\heichips25_can_lehmann_fsm/net916 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1620_  (.Y(\heichips25_can_lehmann_fsm/_0944_ ),
    .A(\heichips25_can_lehmann_fsm/net976 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1621_  (.Y(\heichips25_can_lehmann_fsm/_0945_ ),
    .A(\heichips25_can_lehmann_fsm/net879 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1622_  (.Y(\heichips25_can_lehmann_fsm/_0946_ ),
    .A(\heichips25_can_lehmann_fsm/net1095 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1623_  (.Y(\heichips25_can_lehmann_fsm/_0947_ ),
    .A(\heichips25_can_lehmann_fsm/net1000 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1624_  (.Y(\heichips25_can_lehmann_fsm/_0948_ ),
    .A(\heichips25_can_lehmann_fsm/net1055 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1625_  (.Y(\heichips25_can_lehmann_fsm/_0949_ ),
    .A(\heichips25_can_lehmann_fsm/net1126 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1626_  (.Y(\heichips25_can_lehmann_fsm/_0950_ ),
    .A(\heichips25_can_lehmann_fsm/net1110 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1627_  (.Y(\heichips25_can_lehmann_fsm/_0951_ ),
    .A(\heichips25_can_lehmann_fsm/net1015 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1628_  (.Y(\heichips25_can_lehmann_fsm/_0952_ ),
    .A(\heichips25_can_lehmann_fsm/net1066 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1629_  (.Y(\heichips25_can_lehmann_fsm/_0953_ ),
    .A(\heichips25_can_lehmann_fsm/net1167 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1630_  (.Y(\heichips25_can_lehmann_fsm/_0954_ ),
    .A(\heichips25_can_lehmann_fsm/net987 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1631_  (.Y(\heichips25_can_lehmann_fsm/_0955_ ),
    .A(\heichips25_can_lehmann_fsm/net922 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1632_  (.Y(\heichips25_can_lehmann_fsm/_0956_ ),
    .A(\heichips25_can_lehmann_fsm/net883 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1633_  (.Y(\heichips25_can_lehmann_fsm/_0957_ ),
    .A(\heichips25_can_lehmann_fsm/net1085 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1634_  (.Y(\heichips25_can_lehmann_fsm/_0958_ ),
    .A(\heichips25_can_lehmann_fsm/net948 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1635_  (.Y(\heichips25_can_lehmann_fsm/_0959_ ),
    .A(\heichips25_can_lehmann_fsm/net942 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1636_  (.Y(\heichips25_can_lehmann_fsm/_0960_ ),
    .A(\heichips25_can_lehmann_fsm/net965 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1637_  (.Y(\heichips25_can_lehmann_fsm/_0961_ ),
    .A(\heichips25_can_lehmann_fsm/net939 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1638_  (.Y(\heichips25_can_lehmann_fsm/_0962_ ),
    .A(\heichips25_can_lehmann_fsm/net898 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1639_  (.Y(\heichips25_can_lehmann_fsm/_0963_ ),
    .A(\heichips25_can_lehmann_fsm/net840 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1640_  (.Y(\heichips25_can_lehmann_fsm/_0964_ ),
    .A(\heichips25_can_lehmann_fsm/net1002 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1641_  (.Y(\heichips25_can_lehmann_fsm/_0965_ ),
    .A(\heichips25_can_lehmann_fsm/net1050 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1642_  (.Y(\heichips25_can_lehmann_fsm/_0966_ ),
    .A(\heichips25_can_lehmann_fsm/net1006 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1643_  (.Y(\heichips25_can_lehmann_fsm/_0967_ ),
    .A(\heichips25_can_lehmann_fsm/net851 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1644_  (.Y(\heichips25_can_lehmann_fsm/_0968_ ),
    .A(\heichips25_can_lehmann_fsm/net1088 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1645_  (.Y(\heichips25_can_lehmann_fsm/_0969_ ),
    .A(\heichips25_can_lehmann_fsm/net1099 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1646_  (.Y(\heichips25_can_lehmann_fsm/_0970_ ),
    .A(\heichips25_can_lehmann_fsm/net895 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1647_  (.Y(\heichips25_can_lehmann_fsm/_0971_ ),
    .A(\heichips25_can_lehmann_fsm/net1093 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1648_  (.Y(\heichips25_can_lehmann_fsm/_0972_ ),
    .A(net11));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1649_  (.Y(\heichips25_can_lehmann_fsm/_0973_ ),
    .A(\heichips25_can_lehmann_fsm/net1182 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1650_  (.Y(\heichips25_can_lehmann_fsm/_0974_ ),
    .A(\heichips25_can_lehmann_fsm/net1198 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1651_  (.Y(\heichips25_can_lehmann_fsm/_0975_ ),
    .A(\heichips25_can_lehmann_fsm/net1226 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1652_  (.Y(\heichips25_can_lehmann_fsm/_0976_ ),
    .A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[3] ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1653_  (.Y(\heichips25_can_lehmann_fsm/_0977_ ),
    .A(\heichips25_can_lehmann_fsm/net1255 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1654_  (.Y(\heichips25_can_lehmann_fsm/_0978_ ),
    .A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[23] ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1655_  (.Y(\heichips25_can_lehmann_fsm/_0979_ ),
    .A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[22] ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1656_  (.Y(\heichips25_can_lehmann_fsm/_0980_ ),
    .A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[21] ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1657_  (.Y(\heichips25_can_lehmann_fsm/_0981_ ),
    .A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[16] ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1658_  (.Y(\heichips25_can_lehmann_fsm/_0982_ ),
    .A(\heichips25_can_lehmann_fsm/net1234 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1659_  (.Y(\heichips25_can_lehmann_fsm/_0983_ ),
    .A(\heichips25_can_lehmann_fsm/net348 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1660_  (.Y(\heichips25_can_lehmann_fsm/_0984_ ),
    .A(\heichips25_can_lehmann_fsm/net353 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1661_  (.Y(\heichips25_can_lehmann_fsm/_0985_ ),
    .A(net3));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1662_  (.Y(\heichips25_can_lehmann_fsm/_0986_ ),
    .A(net4));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1663_  (.Y(\heichips25_can_lehmann_fsm/_0987_ ),
    .A(net5));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1664_  (.Y(\heichips25_can_lehmann_fsm/_0988_ ),
    .A(net6));
 sg13g2_nor2b_1 \heichips25_can_lehmann_fsm/_1665_  (.A(\heichips25_can_lehmann_fsm/net351 ),
    .B_N(\heichips25_can_lehmann_fsm/net353 ),
    .Y(\heichips25_can_lehmann_fsm/_0989_ ));
 sg13g2_and2_1 \heichips25_can_lehmann_fsm/_1666_  (.A(\heichips25_can_lehmann_fsm/net350 ),
    .B(\heichips25_can_lehmann_fsm/_0989_ ),
    .X(\heichips25_can_lehmann_fsm/_0990_ ));
 sg13g2_nand3b_1 \heichips25_can_lehmann_fsm/_1667_  (.B(\heichips25_can_lehmann_fsm/net353 ),
    .C(\heichips25_can_lehmann_fsm/net350 ),
    .Y(\heichips25_can_lehmann_fsm/_0991_ ),
    .A_N(\heichips25_can_lehmann_fsm/net351 ));
 sg13g2_nor2b_1 \heichips25_can_lehmann_fsm/_1668_  (.A(\heichips25_can_lehmann_fsm/net353 ),
    .B_N(\heichips25_can_lehmann_fsm/net351 ),
    .Y(\heichips25_can_lehmann_fsm/_0992_ ));
 sg13g2_and2_1 \heichips25_can_lehmann_fsm/_1669_  (.A(\heichips25_can_lehmann_fsm/net338 ),
    .B(\heichips25_can_lehmann_fsm/_0992_ ),
    .X(\heichips25_can_lehmann_fsm/_0993_ ));
 sg13g2_and2_1 \heichips25_can_lehmann_fsm/_1670_  (.A(\heichips25_can_lehmann_fsm/net350 ),
    .B(\heichips25_can_lehmann_fsm/_0992_ ),
    .X(\heichips25_can_lehmann_fsm/_0994_ ));
 sg13g2_nand3b_1 \heichips25_can_lehmann_fsm/_1671_  (.B(\heichips25_can_lehmann_fsm/net351 ),
    .C(\heichips25_can_lehmann_fsm/net348 ),
    .Y(\heichips25_can_lehmann_fsm/_0995_ ),
    .A_N(\heichips25_can_lehmann_fsm/net353 ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_1672_  (.Y(\heichips25_can_lehmann_fsm/_0996_ ),
    .A(\heichips25_can_lehmann_fsm/net352 ),
    .B(\heichips25_can_lehmann_fsm/net353 ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_1673_  (.A(\heichips25_can_lehmann_fsm/net348 ),
    .B(\heichips25_can_lehmann_fsm/_0996_ ),
    .Y(\heichips25_can_lehmann_fsm/_0997_ ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_1674_  (.A(\heichips25_can_lehmann_fsm/net352 ),
    .B(\heichips25_can_lehmann_fsm/net353 ),
    .Y(\heichips25_can_lehmann_fsm/_0998_ ));
 sg13g2_or2_1 \heichips25_can_lehmann_fsm/_1675_  (.X(\heichips25_can_lehmann_fsm/_0999_ ),
    .B(\heichips25_can_lehmann_fsm/net353 ),
    .A(\heichips25_can_lehmann_fsm/net352 ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_1676_  (.A(\heichips25_can_lehmann_fsm/net348 ),
    .B(\heichips25_can_lehmann_fsm/_0999_ ),
    .Y(\heichips25_can_lehmann_fsm/_1000_ ));
 sg13g2_or3_1 \heichips25_can_lehmann_fsm/_1677_  (.A(\heichips25_can_lehmann_fsm/net350 ),
    .B(\heichips25_can_lehmann_fsm/net351 ),
    .C(\heichips25_can_lehmann_fsm/net354 ),
    .X(\heichips25_can_lehmann_fsm/_1001_ ));
 sg13g2_and2_1 \heichips25_can_lehmann_fsm/_1678_  (.A(\heichips25_can_lehmann_fsm/net338 ),
    .B(\heichips25_can_lehmann_fsm/_0989_ ),
    .X(\heichips25_can_lehmann_fsm/_1002_ ));
 sg13g2_and3_1 \heichips25_can_lehmann_fsm/_1679_  (.X(\heichips25_can_lehmann_fsm/_1003_ ),
    .A(\heichips25_can_lehmann_fsm/net350 ),
    .B(\heichips25_can_lehmann_fsm/net351 ),
    .C(\heichips25_can_lehmann_fsm/net354 ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_1680_  (.A(\heichips25_can_lehmann_fsm/net338 ),
    .B(\heichips25_can_lehmann_fsm/_0999_ ),
    .Y(\heichips25_can_lehmann_fsm/_1004_ ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1681_  (.Y(\heichips25_can_lehmann_fsm/_1005_ ),
    .B1(\heichips25_can_lehmann_fsm/net296 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[63] ),
    .A2(\heichips25_can_lehmann_fsm/net317 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[159] ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1682_  (.Y(\heichips25_can_lehmann_fsm/_1006_ ),
    .B1(\heichips25_can_lehmann_fsm/net294 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[135] ),
    .A2(\heichips25_can_lehmann_fsm/net310 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[183] ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1683_  (.Y(\heichips25_can_lehmann_fsm/_1007_ ),
    .B1(\heichips25_can_lehmann_fsm/net331 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[7] ),
    .A2(\heichips25_can_lehmann_fsm/net313 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[87] ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_1684_  (.A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[111] ),
    .A2(\heichips25_can_lehmann_fsm/net305 ),
    .Y(\heichips25_can_lehmann_fsm/_1008_ ),
    .B1(\heichips25_can_lehmann_fsm/net300 ));
 sg13g2_nand4_1 \heichips25_can_lehmann_fsm/_1685_  (.B(\heichips25_can_lehmann_fsm/_1006_ ),
    .C(\heichips25_can_lehmann_fsm/_1007_ ),
    .A(\heichips25_can_lehmann_fsm/_1005_ ),
    .Y(\heichips25_can_lehmann_fsm/_1009_ ),
    .D(\heichips25_can_lehmann_fsm/_1008_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_1686_  (.B1(\heichips25_can_lehmann_fsm/_1009_ ),
    .Y(\heichips25_can_lehmann_fsm/_1010_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[39] ),
    .A2(\heichips25_can_lehmann_fsm/net336 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_1687_  (.A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[112] ),
    .A2(\heichips25_can_lehmann_fsm/net305 ),
    .Y(\heichips25_can_lehmann_fsm/_1011_ ),
    .B1(\heichips25_can_lehmann_fsm/net300 ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1688_  (.Y(\heichips25_can_lehmann_fsm/_1012_ ),
    .B1(\heichips25_can_lehmann_fsm/net296 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[64] ),
    .A2(\heichips25_can_lehmann_fsm/net317 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[160] ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1689_  (.Y(\heichips25_can_lehmann_fsm/_1013_ ),
    .B1(\heichips25_can_lehmann_fsm/net294 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[136] ),
    .A2(\heichips25_can_lehmann_fsm/net310 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[184] ));
 sg13g2_nand3_1 \heichips25_can_lehmann_fsm/_1690_  (.B(\heichips25_can_lehmann_fsm/_1012_ ),
    .C(\heichips25_can_lehmann_fsm/_1013_ ),
    .A(\heichips25_can_lehmann_fsm/_1011_ ),
    .Y(\heichips25_can_lehmann_fsm/_1014_ ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_1691_  (.B2(\heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[8] ),
    .C1(\heichips25_can_lehmann_fsm/_1014_ ),
    .B1(\heichips25_can_lehmann_fsm/net331 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[88] ),
    .Y(\heichips25_can_lehmann_fsm/_1015_ ),
    .A2(\heichips25_can_lehmann_fsm/net313 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_1692_  (.A1(\heichips25_can_lehmann_fsm/_0951_ ),
    .A2(\heichips25_can_lehmann_fsm/net300 ),
    .Y(\heichips25_can_lehmann_fsm/_1016_ ),
    .B1(\heichips25_can_lehmann_fsm/_1015_ ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1693_  (.Y(\heichips25_can_lehmann_fsm/_1017_ ),
    .B1(\heichips25_can_lehmann_fsm/net294 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[134] ),
    .A2(\heichips25_can_lehmann_fsm/net331 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[6] ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1694_  (.Y(\heichips25_can_lehmann_fsm/_1018_ ),
    .B1(\heichips25_can_lehmann_fsm/net296 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[62] ),
    .A2(\heichips25_can_lehmann_fsm/net317 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[158] ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1695_  (.Y(\heichips25_can_lehmann_fsm/_1019_ ),
    .B1(\heichips25_can_lehmann_fsm/net305 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[110] ),
    .A2(\heichips25_can_lehmann_fsm/net313 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[86] ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_1696_  (.A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[182] ),
    .A2(\heichips25_can_lehmann_fsm/net310 ),
    .Y(\heichips25_can_lehmann_fsm/_1020_ ),
    .B1(\heichips25_can_lehmann_fsm/net300 ));
 sg13g2_nand4_1 \heichips25_can_lehmann_fsm/_1697_  (.B(\heichips25_can_lehmann_fsm/_1018_ ),
    .C(\heichips25_can_lehmann_fsm/_1019_ ),
    .A(\heichips25_can_lehmann_fsm/_1017_ ),
    .Y(\heichips25_can_lehmann_fsm/_1021_ ),
    .D(\heichips25_can_lehmann_fsm/_1020_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_1698_  (.B1(\heichips25_can_lehmann_fsm/_1021_ ),
    .Y(\heichips25_can_lehmann_fsm/_1022_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[38] ),
    .A2(\heichips25_can_lehmann_fsm/net336 ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1699_  (.Y(\heichips25_can_lehmann_fsm/_1023_ ),
    .B1(\heichips25_can_lehmann_fsm/net294 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[133] ),
    .A2(\heichips25_can_lehmann_fsm/net317 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[157] ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1700_  (.Y(\heichips25_can_lehmann_fsm/_1024_ ),
    .B1(\heichips25_can_lehmann_fsm/net296 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[61] ),
    .A2(\heichips25_can_lehmann_fsm/net313 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[85] ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_1701_  (.A1(\heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[5] ),
    .A2(\heichips25_can_lehmann_fsm/net331 ),
    .Y(\heichips25_can_lehmann_fsm/_1025_ ),
    .B1(\heichips25_can_lehmann_fsm/net300 ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_1702_  (.Y(\heichips25_can_lehmann_fsm/_1026_ ),
    .A(\heichips25_can_lehmann_fsm/_1024_ ),
    .B(\heichips25_can_lehmann_fsm/_1025_ ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_1703_  (.B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[109] ),
    .C1(\heichips25_can_lehmann_fsm/_1026_ ),
    .B1(\heichips25_can_lehmann_fsm/net305 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[181] ),
    .Y(\heichips25_can_lehmann_fsm/_1027_ ),
    .A2(\heichips25_can_lehmann_fsm/net310 ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1704_  (.Y(\heichips25_can_lehmann_fsm/_1028_ ),
    .B1(\heichips25_can_lehmann_fsm/_1023_ ),
    .B2(\heichips25_can_lehmann_fsm/_1027_ ),
    .A2(\heichips25_can_lehmann_fsm/net300 ),
    .A1(\heichips25_can_lehmann_fsm/_0953_ ));
 sg13g2_nand2b_1 \heichips25_can_lehmann_fsm/_1705_  (.Y(\heichips25_can_lehmann_fsm/_1029_ ),
    .B(\heichips25_can_lehmann_fsm/_1028_ ),
    .A_N(\heichips25_can_lehmann_fsm/_1022_ ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_1706_  (.A(\heichips25_can_lehmann_fsm/_1016_ ),
    .B(\heichips25_can_lehmann_fsm/_1029_ ),
    .Y(\heichips25_can_lehmann_fsm/_1030_ ));
 sg13g2_or2_1 \heichips25_can_lehmann_fsm/_1707_  (.X(\heichips25_can_lehmann_fsm/_1031_ ),
    .B(\heichips25_can_lehmann_fsm/_1029_ ),
    .A(\heichips25_can_lehmann_fsm/_1016_ ));
 sg13g2_and2_1 \heichips25_can_lehmann_fsm/_1708_  (.A(\heichips25_can_lehmann_fsm/_1010_ ),
    .B(\heichips25_can_lehmann_fsm/_1030_ ),
    .X(\heichips25_can_lehmann_fsm/_1032_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_1709_  (.A1(\heichips25_can_lehmann_fsm/_1022_ ),
    .A2(\heichips25_can_lehmann_fsm/_1028_ ),
    .Y(\heichips25_can_lehmann_fsm/_1033_ ),
    .B1(\heichips25_can_lehmann_fsm/_1032_ ));
 sg13g2_nor2b_1 \heichips25_can_lehmann_fsm/_1710_  (.A(\heichips25_can_lehmann_fsm/_1010_ ),
    .B_N(\heichips25_can_lehmann_fsm/_1016_ ),
    .Y(\heichips25_can_lehmann_fsm/_1034_ ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_1711_  (.Y(\heichips25_can_lehmann_fsm/_1035_ ),
    .A(\heichips25_can_lehmann_fsm/controller.output_controller.keep[0] ),
    .B(\heichips25_can_lehmann_fsm/_1034_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_1712_  (.A1(\heichips25_can_lehmann_fsm/_1028_ ),
    .A2(\heichips25_can_lehmann_fsm/_1035_ ),
    .Y(\heichips25_can_lehmann_fsm/_1036_ ),
    .B1(\heichips25_can_lehmann_fsm/_1022_ ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_1713_  (.A(\heichips25_can_lehmann_fsm/_1010_ ),
    .B(\heichips25_can_lehmann_fsm/_1031_ ),
    .Y(\heichips25_can_lehmann_fsm/_1037_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_1714_  (.A1(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[16] ),
    .A2(\heichips25_can_lehmann_fsm/_1037_ ),
    .Y(\heichips25_can_lehmann_fsm/_1038_ ),
    .B1(\heichips25_can_lehmann_fsm/_1036_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_1715_  (.B1(\heichips25_can_lehmann_fsm/_1038_ ),
    .Y(\uo_out_fsm[0] ),
    .A1(\heichips25_can_lehmann_fsm/_0977_ ),
    .A2(\heichips25_can_lehmann_fsm/_1033_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_1716_  (.A1(\heichips25_can_lehmann_fsm/net1277 ),
    .A2(\heichips25_can_lehmann_fsm/_1016_ ),
    .Y(\heichips25_can_lehmann_fsm/_1039_ ),
    .B1(\heichips25_can_lehmann_fsm/_1029_ ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1717_  (.Y(\heichips25_can_lehmann_fsm/_1040_ ),
    .B1(\heichips25_can_lehmann_fsm/_1037_ ),
    .B2(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[17] ),
    .A2(\heichips25_can_lehmann_fsm/_1032_ ),
    .A1(\heichips25_can_lehmann_fsm/net347 ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_1718_  (.B1(\heichips25_can_lehmann_fsm/_1040_ ),
    .Y(\uo_out_fsm[1] ),
    .A1(\heichips25_can_lehmann_fsm/_1010_ ),
    .A2(\heichips25_can_lehmann_fsm/_1039_ ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1719_  (.Y(\heichips25_can_lehmann_fsm/_1041_ ),
    .B1(\heichips25_can_lehmann_fsm/_1034_ ),
    .B2(\heichips25_can_lehmann_fsm/net1213 ),
    .A2(\heichips25_can_lehmann_fsm/_1029_ ),
    .A1(\heichips25_can_lehmann_fsm/_1016_ ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1720_  (.Y(\heichips25_can_lehmann_fsm/_1042_ ),
    .B1(\heichips25_can_lehmann_fsm/_1037_ ),
    .B2(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[18] ),
    .A2(\heichips25_can_lehmann_fsm/_1032_ ),
    .A1(\heichips25_can_lehmann_fsm/net346 ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_1721_  (.Y(\uo_out_fsm[2] ),
    .A(\heichips25_can_lehmann_fsm/_1041_ ),
    .B(\heichips25_can_lehmann_fsm/_1042_ ));
 sg13g2_nor3_1 \heichips25_can_lehmann_fsm/_1722_  (.A(\heichips25_can_lehmann_fsm/net1195 ),
    .B(\heichips25_can_lehmann_fsm/net1174 ),
    .C(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[0] ),
    .Y(\heichips25_can_lehmann_fsm/_1043_ ));
 sg13g2_or4_1 \heichips25_can_lehmann_fsm/_1723_  (.A(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[3] ),
    .B(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[2] ),
    .C(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[1] ),
    .D(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[0] ),
    .X(\heichips25_can_lehmann_fsm/_1044_ ));
 sg13g2_nor3_1 \heichips25_can_lehmann_fsm/_1724_  (.A(\heichips25_can_lehmann_fsm/net1181 ),
    .B(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[4] ),
    .C(\heichips25_can_lehmann_fsm/_1044_ ),
    .Y(\heichips25_can_lehmann_fsm/_1045_ ));
 sg13g2_nor4_1 \heichips25_can_lehmann_fsm/_1725_  (.A(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[6] ),
    .B(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[5] ),
    .C(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[4] ),
    .D(\heichips25_can_lehmann_fsm/_1044_ ),
    .Y(\heichips25_can_lehmann_fsm/_1046_ ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_1726_  (.Y(\heichips25_can_lehmann_fsm/_1047_ ),
    .A(\heichips25_can_lehmann_fsm/_0973_ ),
    .B(\heichips25_can_lehmann_fsm/_1046_ ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_1727_  (.A(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[9] ),
    .B(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[8] ),
    .Y(\heichips25_can_lehmann_fsm/_1048_ ));
 sg13g2_nand3_1 \heichips25_can_lehmann_fsm/_1728_  (.B(\heichips25_can_lehmann_fsm/_1046_ ),
    .C(\heichips25_can_lehmann_fsm/_1048_ ),
    .A(\heichips25_can_lehmann_fsm/_0973_ ),
    .Y(\heichips25_can_lehmann_fsm/_1049_ ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_1729_  (.A(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[11] ),
    .B(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[10] ),
    .Y(\heichips25_can_lehmann_fsm/_1050_ ));
 sg13g2_nand4_1 \heichips25_can_lehmann_fsm/_1730_  (.B(\heichips25_can_lehmann_fsm/_1046_ ),
    .C(\heichips25_can_lehmann_fsm/_1048_ ),
    .A(\heichips25_can_lehmann_fsm/_0973_ ),
    .Y(\heichips25_can_lehmann_fsm/_1051_ ),
    .D(\heichips25_can_lehmann_fsm/_1050_ ));
 sg13g2_nor3_1 \heichips25_can_lehmann_fsm/_1731_  (.A(\heichips25_can_lehmann_fsm/net1158 ),
    .B(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[12] ),
    .C(\heichips25_can_lehmann_fsm/_1051_ ),
    .Y(\heichips25_can_lehmann_fsm/_1052_ ));
 sg13g2_nor4_1 \heichips25_can_lehmann_fsm/_1732_  (.A(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[15] ),
    .B(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[14] ),
    .C(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[13] ),
    .D(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[12] ),
    .Y(\heichips25_can_lehmann_fsm/_1053_ ));
 sg13g2_nand2b_1 \heichips25_can_lehmann_fsm/_1733_  (.Y(\heichips25_can_lehmann_fsm/_1054_ ),
    .B(\heichips25_can_lehmann_fsm/_1053_ ),
    .A_N(\heichips25_can_lehmann_fsm/_1051_ ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1734_  (.Y(\heichips25_can_lehmann_fsm/_1055_ ),
    .B1(\heichips25_can_lehmann_fsm/_1037_ ),
    .B2(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[19] ),
    .A2(\heichips25_can_lehmann_fsm/_1032_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[3] ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_1735_  (.B1(\heichips25_can_lehmann_fsm/_1055_ ),
    .Y(\uo_out_fsm[3] ),
    .A1(\heichips25_can_lehmann_fsm/_1030_ ),
    .A2(\heichips25_can_lehmann_fsm/_1054_ ));
 sg13g2_or4_1 \heichips25_can_lehmann_fsm/_1736_  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[3] ),
    .B(\heichips25_can_lehmann_fsm/net346 ),
    .C(\heichips25_can_lehmann_fsm/net347 ),
    .D(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[0] ),
    .X(\heichips25_can_lehmann_fsm/_1056_ ));
 sg13g2_or2_1 \heichips25_can_lehmann_fsm/_1737_  (.X(\heichips25_can_lehmann_fsm/_1057_ ),
    .B(\heichips25_can_lehmann_fsm/net345 ),
    .A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[5] ));
 sg13g2_or2_1 \heichips25_can_lehmann_fsm/_1738_  (.X(\heichips25_can_lehmann_fsm/_1058_ ),
    .B(\heichips25_can_lehmann_fsm/_1057_ ),
    .A(\heichips25_can_lehmann_fsm/_1056_ ));
 sg13g2_or2_1 \heichips25_can_lehmann_fsm/_1739_  (.X(\heichips25_can_lehmann_fsm/_1059_ ),
    .B(\heichips25_can_lehmann_fsm/net344 ),
    .A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[7] ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_1740_  (.A(\heichips25_can_lehmann_fsm/_1058_ ),
    .B(\heichips25_can_lehmann_fsm/_1059_ ),
    .Y(\heichips25_can_lehmann_fsm/_1060_ ));
 sg13g2_nor4_1 \heichips25_can_lehmann_fsm/_1741_  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[8] ),
    .B(\heichips25_can_lehmann_fsm/_1056_ ),
    .C(\heichips25_can_lehmann_fsm/_1057_ ),
    .D(\heichips25_can_lehmann_fsm/_1059_ ),
    .Y(\heichips25_can_lehmann_fsm/_1061_ ));
 sg13g2_nor2b_1 \heichips25_can_lehmann_fsm/_1742_  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[9] ),
    .B_N(\heichips25_can_lehmann_fsm/_1061_ ),
    .Y(\heichips25_can_lehmann_fsm/_1062_ ));
 sg13g2_nand2b_1 \heichips25_can_lehmann_fsm/_1743_  (.Y(\heichips25_can_lehmann_fsm/_1063_ ),
    .B(\heichips25_can_lehmann_fsm/_1062_ ),
    .A_N(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[10] ));
 sg13g2_nor3_1 \heichips25_can_lehmann_fsm/_1744_  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[11] ),
    .B(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[10] ),
    .C(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[9] ),
    .Y(\heichips25_can_lehmann_fsm/_1064_ ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_1745_  (.Y(\heichips25_can_lehmann_fsm/_1065_ ),
    .A(\heichips25_can_lehmann_fsm/_1061_ ),
    .B(\heichips25_can_lehmann_fsm/_1064_ ));
 sg13g2_nor4_1 \heichips25_can_lehmann_fsm/_1746_  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[15] ),
    .B(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[14] ),
    .C(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[13] ),
    .D(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[12] ),
    .Y(\heichips25_can_lehmann_fsm/_1066_ ));
 sg13g2_nand3_1 \heichips25_can_lehmann_fsm/_1747_  (.B(\heichips25_can_lehmann_fsm/_1064_ ),
    .C(\heichips25_can_lehmann_fsm/_1066_ ),
    .A(\heichips25_can_lehmann_fsm/_1061_ ),
    .Y(\heichips25_can_lehmann_fsm/_1067_ ));
 sg13g2_nand4_1 \heichips25_can_lehmann_fsm/_1748_  (.B(\heichips25_can_lehmann_fsm/_1061_ ),
    .C(\heichips25_can_lehmann_fsm/_1064_ ),
    .A(\heichips25_can_lehmann_fsm/_0981_ ),
    .Y(\heichips25_can_lehmann_fsm/_1068_ ),
    .D(\heichips25_can_lehmann_fsm/_1066_ ));
 sg13g2_or2_1 \heichips25_can_lehmann_fsm/_1749_  (.X(\heichips25_can_lehmann_fsm/_1069_ ),
    .B(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[17] ),
    .A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[18] ));
 sg13g2_or2_1 \heichips25_can_lehmann_fsm/_1750_  (.X(\heichips25_can_lehmann_fsm/_1070_ ),
    .B(\heichips25_can_lehmann_fsm/_1069_ ),
    .A(\heichips25_can_lehmann_fsm/_1068_ ));
 sg13g2_nor4_1 \heichips25_can_lehmann_fsm/_1751_  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[20] ),
    .B(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[19] ),
    .C(\heichips25_can_lehmann_fsm/_1068_ ),
    .D(\heichips25_can_lehmann_fsm/_1069_ ),
    .Y(\heichips25_can_lehmann_fsm/_1071_ ));
 sg13g2_or4_1 \heichips25_can_lehmann_fsm/_1752_  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[20] ),
    .B(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[19] ),
    .C(\heichips25_can_lehmann_fsm/_1068_ ),
    .D(\heichips25_can_lehmann_fsm/_1069_ ),
    .X(\heichips25_can_lehmann_fsm/_1072_ ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_1753_  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[21] ),
    .B(\heichips25_can_lehmann_fsm/_1072_ ),
    .Y(\heichips25_can_lehmann_fsm/_1073_ ));
 sg13g2_nor4_1 \heichips25_can_lehmann_fsm/_1754_  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[23] ),
    .B(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[22] ),
    .C(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[21] ),
    .D(\heichips25_can_lehmann_fsm/_1072_ ),
    .Y(\heichips25_can_lehmann_fsm/_1074_ ));
 sg13g2_nand4_1 \heichips25_can_lehmann_fsm/_1755_  (.B(\heichips25_can_lehmann_fsm/_0979_ ),
    .C(\heichips25_can_lehmann_fsm/_0980_ ),
    .A(\heichips25_can_lehmann_fsm/_0978_ ),
    .Y(\heichips25_can_lehmann_fsm/_1075_ ),
    .D(\heichips25_can_lehmann_fsm/_1071_ ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_1756_  (.Y(\heichips25_can_lehmann_fsm/_1076_ ),
    .A(\heichips25_can_lehmann_fsm/net345 ),
    .B(\heichips25_can_lehmann_fsm/_1032_ ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1757_  (.Y(\heichips25_can_lehmann_fsm/_1077_ ),
    .B1(\heichips25_can_lehmann_fsm/_1074_ ),
    .B2(\heichips25_can_lehmann_fsm/_1031_ ),
    .A2(\heichips25_can_lehmann_fsm/_1037_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[20] ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_1758_  (.Y(\uo_out_fsm[4] ),
    .A(\heichips25_can_lehmann_fsm/_1076_ ),
    .B(\heichips25_can_lehmann_fsm/_1077_ ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_1759_  (.Y(\heichips25_can_lehmann_fsm/_1078_ ),
    .A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[21] ),
    .B(\heichips25_can_lehmann_fsm/_1037_ ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1760_  (.Y(\heichips25_can_lehmann_fsm/_1079_ ),
    .B1(\heichips25_can_lehmann_fsm/_1032_ ),
    .B2(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[5] ),
    .A2(\heichips25_can_lehmann_fsm/_1031_ ),
    .A1(\heichips25_can_lehmann_fsm/net354 ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_1761_  (.Y(\uo_out_fsm[5] ),
    .A(\heichips25_can_lehmann_fsm/_1078_ ),
    .B(\heichips25_can_lehmann_fsm/_1079_ ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_1762_  (.Y(\heichips25_can_lehmann_fsm/_1080_ ),
    .A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[22] ),
    .B(\heichips25_can_lehmann_fsm/_1037_ ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1763_  (.Y(\heichips25_can_lehmann_fsm/_1081_ ),
    .B1(\heichips25_can_lehmann_fsm/_1032_ ),
    .B2(\heichips25_can_lehmann_fsm/net344 ),
    .A2(\heichips25_can_lehmann_fsm/_1031_ ),
    .A1(\heichips25_can_lehmann_fsm/net351 ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_1764_  (.Y(\uo_out_fsm[6] ),
    .A(\heichips25_can_lehmann_fsm/_1080_ ),
    .B(\heichips25_can_lehmann_fsm/_1081_ ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_1765_  (.Y(\heichips25_can_lehmann_fsm/_1082_ ),
    .A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[23] ),
    .B(\heichips25_can_lehmann_fsm/_1037_ ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1766_  (.Y(\heichips25_can_lehmann_fsm/_1083_ ),
    .B1(\heichips25_can_lehmann_fsm/_1032_ ),
    .B2(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[7] ),
    .A2(\heichips25_can_lehmann_fsm/_1031_ ),
    .A1(\heichips25_can_lehmann_fsm/net350 ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_1767_  (.Y(\uo_out_fsm[7] ),
    .A(\heichips25_can_lehmann_fsm/_1082_ ),
    .B(\heichips25_can_lehmann_fsm/_1083_ ));
 sg13g2_or2_1 \heichips25_can_lehmann_fsm/_1768_  (.X(\heichips25_can_lehmann_fsm/_1084_ ),
    .B(\heichips25_can_lehmann_fsm/net335 ),
    .A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[36] ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1769_  (.Y(\heichips25_can_lehmann_fsm/_1085_ ),
    .B1(\heichips25_can_lehmann_fsm/net331 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[4] ),
    .A2(\heichips25_can_lehmann_fsm/net317 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[156] ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1770_  (.Y(\heichips25_can_lehmann_fsm/_1086_ ),
    .B1(\heichips25_can_lehmann_fsm/net310 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[180] ),
    .A2(\heichips25_can_lehmann_fsm/net313 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[84] ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1771_  (.Y(\heichips25_can_lehmann_fsm/_1087_ ),
    .B1(\heichips25_can_lehmann_fsm/net294 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[132] ),
    .A2(\heichips25_can_lehmann_fsm/net305 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[108] ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_1772_  (.A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[60] ),
    .A2(\heichips25_can_lehmann_fsm/net296 ),
    .Y(\heichips25_can_lehmann_fsm/_1088_ ),
    .B1(\heichips25_can_lehmann_fsm/net300 ));
 sg13g2_nand4_1 \heichips25_can_lehmann_fsm/_1773_  (.B(\heichips25_can_lehmann_fsm/_1086_ ),
    .C(\heichips25_can_lehmann_fsm/_1087_ ),
    .A(\heichips25_can_lehmann_fsm/_1085_ ),
    .Y(\heichips25_can_lehmann_fsm/_1089_ ),
    .D(\heichips25_can_lehmann_fsm/_1088_ ));
 sg13g2_nand3_1 \heichips25_can_lehmann_fsm/_1774_  (.B(\heichips25_can_lehmann_fsm/_1084_ ),
    .C(\heichips25_can_lehmann_fsm/_1089_ ),
    .A(\heichips25_can_lehmann_fsm/_1054_ ),
    .Y(\heichips25_can_lehmann_fsm/_1090_ ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1775_  (.Y(\heichips25_can_lehmann_fsm/_1091_ ),
    .B1(\heichips25_can_lehmann_fsm/net332 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[3] ),
    .A2(\heichips25_can_lehmann_fsm/net317 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[155] ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1776_  (.Y(\heichips25_can_lehmann_fsm/_1092_ ),
    .B1(\heichips25_can_lehmann_fsm/net295 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[131] ),
    .A2(\heichips25_can_lehmann_fsm/net296 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[59] ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1777_  (.Y(\heichips25_can_lehmann_fsm/_1093_ ),
    .B1(\heichips25_can_lehmann_fsm/net305 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[107] ),
    .A2(\heichips25_can_lehmann_fsm/net314 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[83] ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_1778_  (.A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[179] ),
    .A2(\heichips25_can_lehmann_fsm/net310 ),
    .Y(\heichips25_can_lehmann_fsm/_1094_ ),
    .B1(\heichips25_can_lehmann_fsm/net302 ));
 sg13g2_nand4_1 \heichips25_can_lehmann_fsm/_1779_  (.B(\heichips25_can_lehmann_fsm/_1092_ ),
    .C(\heichips25_can_lehmann_fsm/_1093_ ),
    .A(\heichips25_can_lehmann_fsm/_1091_ ),
    .Y(\heichips25_can_lehmann_fsm/_1095_ ),
    .D(\heichips25_can_lehmann_fsm/_1094_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_1780_  (.B1(\heichips25_can_lehmann_fsm/_1095_ ),
    .Y(\heichips25_can_lehmann_fsm/_1096_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[35] ),
    .A2(\heichips25_can_lehmann_fsm/net335 ));
 sg13g2_nor3_1 \heichips25_can_lehmann_fsm/_1781_  (.A(\heichips25_can_lehmann_fsm/net1215 ),
    .B(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[1] ),
    .C(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[0] ),
    .Y(\heichips25_can_lehmann_fsm/_1097_ ));
 sg13g2_or4_1 \heichips25_can_lehmann_fsm/_1782_  (.A(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[3] ),
    .B(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[2] ),
    .C(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[1] ),
    .D(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[0] ),
    .X(\heichips25_can_lehmann_fsm/_1098_ ));
 sg13g2_nor3_1 \heichips25_can_lehmann_fsm/_1783_  (.A(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[5] ),
    .B(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[4] ),
    .C(\heichips25_can_lehmann_fsm/_1098_ ),
    .Y(\heichips25_can_lehmann_fsm/_1099_ ));
 sg13g2_nor4_1 \heichips25_can_lehmann_fsm/_1784_  (.A(\heichips25_can_lehmann_fsm/net1192 ),
    .B(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[5] ),
    .C(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[4] ),
    .D(\heichips25_can_lehmann_fsm/_1098_ ),
    .Y(\heichips25_can_lehmann_fsm/_1100_ ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_1785_  (.Y(\heichips25_can_lehmann_fsm/_1101_ ),
    .A(\heichips25_can_lehmann_fsm/_0974_ ),
    .B(\heichips25_can_lehmann_fsm/_1100_ ));
 sg13g2_nand3b_1 \heichips25_can_lehmann_fsm/_1786_  (.B(\heichips25_can_lehmann_fsm/_0974_ ),
    .C(\heichips25_can_lehmann_fsm/_1100_ ),
    .Y(\heichips25_can_lehmann_fsm/_1102_ ),
    .A_N(\heichips25_can_lehmann_fsm/net1278 ));
 sg13g2_or3_1 \heichips25_can_lehmann_fsm/_1787_  (.A(\heichips25_can_lehmann_fsm/net1207 ),
    .B(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[9] ),
    .C(\heichips25_can_lehmann_fsm/_1102_ ),
    .X(\heichips25_can_lehmann_fsm/_1103_ ));
 sg13g2_or4_1 \heichips25_can_lehmann_fsm/_1788_  (.A(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[11] ),
    .B(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[10] ),
    .C(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[9] ),
    .D(\heichips25_can_lehmann_fsm/_1102_ ),
    .X(\heichips25_can_lehmann_fsm/_1104_ ));
 sg13g2_nor3_1 \heichips25_can_lehmann_fsm/_1789_  (.A(\heichips25_can_lehmann_fsm/net1217 ),
    .B(\heichips25_can_lehmann_fsm/net1279 ),
    .C(\heichips25_can_lehmann_fsm/_1104_ ),
    .Y(\heichips25_can_lehmann_fsm/_1105_ ));
 sg13g2_nor2b_1 \heichips25_can_lehmann_fsm/_1790_  (.A(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[14] ),
    .B_N(\heichips25_can_lehmann_fsm/_1105_ ),
    .Y(\heichips25_can_lehmann_fsm/_1106_ ));
 sg13g2_nor4_1 \heichips25_can_lehmann_fsm/_1791_  (.A(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[15] ),
    .B(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[14] ),
    .C(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[13] ),
    .D(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[12] ),
    .Y(\heichips25_can_lehmann_fsm/_1107_ ));
 sg13g2_nand2b_1 \heichips25_can_lehmann_fsm/_1792_  (.Y(\heichips25_can_lehmann_fsm/_1108_ ),
    .B(\heichips25_can_lehmann_fsm/_1107_ ),
    .A_N(\heichips25_can_lehmann_fsm/_1104_ ));
 sg13g2_nand4_1 \heichips25_can_lehmann_fsm/_1793_  (.B(\heichips25_can_lehmann_fsm/net350 ),
    .C(\heichips25_can_lehmann_fsm/net351 ),
    .A(\heichips25_can_lehmann_fsm/controller.extended_cond.opcode[2] ),
    .Y(\heichips25_can_lehmann_fsm/_1109_ ),
    .D(\heichips25_can_lehmann_fsm/net354 ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_1794_  (.B1(\heichips25_can_lehmann_fsm/_1109_ ),
    .Y(\heichips25_can_lehmann_fsm/_1110_ ),
    .A1(\heichips25_can_lehmann_fsm/_0885_ ),
    .A2(\heichips25_can_lehmann_fsm/_0991_ ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_1795_  (.B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[139] ),
    .C1(\heichips25_can_lehmann_fsm/_1110_ ),
    .B1(\heichips25_can_lehmann_fsm/net294 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[115] ),
    .Y(\heichips25_can_lehmann_fsm/_1111_ ),
    .A2(\heichips25_can_lehmann_fsm/net306 ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_1796_  (.B1(\heichips25_can_lehmann_fsm/net336 ),
    .Y(\heichips25_can_lehmann_fsm/_1112_ ),
    .A1(\heichips25_can_lehmann_fsm/_0872_ ),
    .A2(\heichips25_can_lehmann_fsm/_0995_ ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_1797_  (.B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[67] ),
    .C1(\heichips25_can_lehmann_fsm/_1112_ ),
    .B1(\heichips25_can_lehmann_fsm/net296 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[91] ),
    .Y(\heichips25_can_lehmann_fsm/_1113_ ),
    .A2(\heichips25_can_lehmann_fsm/net313 ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1798_  (.Y(\heichips25_can_lehmann_fsm/_1114_ ),
    .B1(\heichips25_can_lehmann_fsm/_1111_ ),
    .B2(\heichips25_can_lehmann_fsm/_1113_ ),
    .A2(\heichips25_can_lehmann_fsm/net301 ),
    .A1(\heichips25_can_lehmann_fsm/_0949_ ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_1799_  (.A(\heichips25_can_lehmann_fsm/_0886_ ),
    .B(\heichips25_can_lehmann_fsm/_0991_ ),
    .Y(\heichips25_can_lehmann_fsm/_1115_ ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_1800_  (.B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[114] ),
    .C1(\heichips25_can_lehmann_fsm/_1115_ ),
    .B1(\heichips25_can_lehmann_fsm/net306 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[186] ),
    .Y(\heichips25_can_lehmann_fsm/_1116_ ),
    .A2(\heichips25_can_lehmann_fsm/net310 ));
 sg13g2_nand3_1 \heichips25_can_lehmann_fsm/_1801_  (.B(\heichips25_can_lehmann_fsm/net338 ),
    .C(\heichips25_can_lehmann_fsm/_0989_ ),
    .A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[66] ),
    .Y(\heichips25_can_lehmann_fsm/_1117_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_1802_  (.B1(\heichips25_can_lehmann_fsm/net337 ),
    .Y(\heichips25_can_lehmann_fsm/_1118_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[138] ),
    .A2(\heichips25_can_lehmann_fsm/net338 ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_1803_  (.Y(\heichips25_can_lehmann_fsm/_1119_ ),
    .A(\heichips25_can_lehmann_fsm/controller.extended_cond.opcode[1] ),
    .B(\heichips25_can_lehmann_fsm/net331 ));
 sg13g2_nand3_1 \heichips25_can_lehmann_fsm/_1804_  (.B(\heichips25_can_lehmann_fsm/net338 ),
    .C(\heichips25_can_lehmann_fsm/_0992_ ),
    .A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[90] ),
    .Y(\heichips25_can_lehmann_fsm/_1120_ ));
 sg13g2_and4_1 \heichips25_can_lehmann_fsm/_1805_  (.A(\heichips25_can_lehmann_fsm/_1117_ ),
    .B(\heichips25_can_lehmann_fsm/_1118_ ),
    .C(\heichips25_can_lehmann_fsm/_1119_ ),
    .D(\heichips25_can_lehmann_fsm/_1120_ ),
    .X(\heichips25_can_lehmann_fsm/_1121_ ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1806_  (.Y(\heichips25_can_lehmann_fsm/_1122_ ),
    .B1(\heichips25_can_lehmann_fsm/_1116_ ),
    .B2(\heichips25_can_lehmann_fsm/_1121_ ),
    .A2(\heichips25_can_lehmann_fsm/net301 ),
    .A1(\heichips25_can_lehmann_fsm/_0950_ ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_1807_  (.A(\heichips25_can_lehmann_fsm/_1114_ ),
    .B(\heichips25_can_lehmann_fsm/_1122_ ),
    .Y(\heichips25_can_lehmann_fsm/_1123_ ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1808_  (.Y(\heichips25_can_lehmann_fsm/_1124_ ),
    .B1(\heichips25_can_lehmann_fsm/net331 ),
    .B2(\heichips25_can_lehmann_fsm/net343 ),
    .A2(\heichips25_can_lehmann_fsm/net313 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[89] ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_1809_  (.A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[65] ),
    .A2(\heichips25_can_lehmann_fsm/net296 ),
    .Y(\heichips25_can_lehmann_fsm/_1125_ ),
    .B1(\heichips25_can_lehmann_fsm/net300 ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1810_  (.Y(\heichips25_can_lehmann_fsm/_1126_ ),
    .B1(\heichips25_can_lehmann_fsm/net294 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[137] ),
    .A2(\heichips25_can_lehmann_fsm/net317 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[161] ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1811_  (.Y(\heichips25_can_lehmann_fsm/_1127_ ),
    .B1(\heichips25_can_lehmann_fsm/net305 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[113] ),
    .A2(\heichips25_can_lehmann_fsm/net310 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[185] ));
 sg13g2_and3_1 \heichips25_can_lehmann_fsm/_1812_  (.X(\heichips25_can_lehmann_fsm/_1128_ ),
    .A(\heichips25_can_lehmann_fsm/_1125_ ),
    .B(\heichips25_can_lehmann_fsm/_1126_ ),
    .C(\heichips25_can_lehmann_fsm/_1127_ ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_1813_  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[41] ),
    .B(\heichips25_can_lehmann_fsm/net336 ),
    .Y(\heichips25_can_lehmann_fsm/_1129_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_1814_  (.A1(\heichips25_can_lehmann_fsm/_1124_ ),
    .A2(\heichips25_can_lehmann_fsm/_1128_ ),
    .Y(\heichips25_can_lehmann_fsm/_1130_ ),
    .B1(\heichips25_can_lehmann_fsm/_1129_ ));
 sg13g2_a21o_1 \heichips25_can_lehmann_fsm/_1815_  (.A2(\heichips25_can_lehmann_fsm/_1128_ ),
    .A1(\heichips25_can_lehmann_fsm/_1124_ ),
    .B1(\heichips25_can_lehmann_fsm/_1129_ ),
    .X(\heichips25_can_lehmann_fsm/_1131_ ));
 sg13g2_mux2_1 \heichips25_can_lehmann_fsm/_1816_  (.A0(\heichips25_can_lehmann_fsm/_0985_ ),
    .A1(\heichips25_can_lehmann_fsm/_0987_ ),
    .S(\heichips25_can_lehmann_fsm/_1122_ ),
    .X(\heichips25_can_lehmann_fsm/_1132_ ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_1817_  (.B2(\heichips25_can_lehmann_fsm/_1114_ ),
    .C1(\heichips25_can_lehmann_fsm/_1130_ ),
    .B1(\heichips25_can_lehmann_fsm/_1132_ ),
    .A1(\heichips25_can_lehmann_fsm/_1108_ ),
    .Y(\heichips25_can_lehmann_fsm/_1133_ ),
    .A2(\heichips25_can_lehmann_fsm/_1123_ ));
 sg13g2_nor2b_1 \heichips25_can_lehmann_fsm/_1818_  (.A(\heichips25_can_lehmann_fsm/_1114_ ),
    .B_N(\heichips25_can_lehmann_fsm/_1122_ ),
    .Y(\heichips25_can_lehmann_fsm/_1134_ ));
 sg13g2_mux2_1 \heichips25_can_lehmann_fsm/_1819_  (.A0(\heichips25_can_lehmann_fsm/_0986_ ),
    .A1(\heichips25_can_lehmann_fsm/_0988_ ),
    .S(\heichips25_can_lehmann_fsm/_1122_ ),
    .X(\heichips25_can_lehmann_fsm/_1135_ ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_1820_  (.Y(\heichips25_can_lehmann_fsm/_1136_ ),
    .A(\heichips25_can_lehmann_fsm/_1054_ ),
    .B(\heichips25_can_lehmann_fsm/_1123_ ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_1821_  (.B2(\heichips25_can_lehmann_fsm/_1114_ ),
    .C1(\heichips25_can_lehmann_fsm/_1131_ ),
    .B1(\heichips25_can_lehmann_fsm/_1135_ ),
    .A1(\heichips25_can_lehmann_fsm/_1075_ ),
    .Y(\heichips25_can_lehmann_fsm/_1137_ ),
    .A2(\heichips25_can_lehmann_fsm/_1134_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_1822_  (.A1(\heichips25_can_lehmann_fsm/_1136_ ),
    .A2(\heichips25_can_lehmann_fsm/_1137_ ),
    .Y(\heichips25_can_lehmann_fsm/_1138_ ),
    .B1(\heichips25_can_lehmann_fsm/_1133_ ));
 sg13g2_a21o_1 \heichips25_can_lehmann_fsm/_1823_  (.A2(\heichips25_can_lehmann_fsm/_1137_ ),
    .A1(\heichips25_can_lehmann_fsm/_1136_ ),
    .B1(\heichips25_can_lehmann_fsm/_1133_ ),
    .X(\heichips25_can_lehmann_fsm/_1139_ ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_1824_  (.A(\heichips25_can_lehmann_fsm/controller.extended_cond.opcode[2] ),
    .B(\heichips25_can_lehmann_fsm/controller.extended_cond.opcode[1] ),
    .Y(\heichips25_can_lehmann_fsm/_1140_ ));
 sg13g2_nor3_1 \heichips25_can_lehmann_fsm/_1825_  (.A(\heichips25_can_lehmann_fsm/controller.extended_cond.opcode[2] ),
    .B(\heichips25_can_lehmann_fsm/controller.extended_cond.opcode[1] ),
    .C(\heichips25_can_lehmann_fsm/net343 ),
    .Y(\heichips25_can_lehmann_fsm/_1141_ ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1826_  (.Y(\heichips25_can_lehmann_fsm/_1142_ ),
    .A(\heichips25_can_lehmann_fsm/_1141_ ));
 sg13g2_nor2b_1 \heichips25_can_lehmann_fsm/_1827_  (.A(\heichips25_can_lehmann_fsm/controller.extended_cond.opcode[2] ),
    .B_N(\heichips25_can_lehmann_fsm/net343 ),
    .Y(\heichips25_can_lehmann_fsm/_1143_ ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_1828_  (.Y(\heichips25_can_lehmann_fsm/_1144_ ),
    .A(\heichips25_can_lehmann_fsm/controller.extended_cond.opcode[1] ),
    .B(\heichips25_can_lehmann_fsm/_1143_ ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_1829_  (.Y(\heichips25_can_lehmann_fsm/_1145_ ),
    .A(\heichips25_can_lehmann_fsm/net343 ),
    .B(net6));
 sg13g2_nand2b_1 \heichips25_can_lehmann_fsm/_1830_  (.Y(\heichips25_can_lehmann_fsm/_1146_ ),
    .B(net5),
    .A_N(\heichips25_can_lehmann_fsm/net343 ));
 sg13g2_nand4_1 \heichips25_can_lehmann_fsm/_1831_  (.B(\heichips25_can_lehmann_fsm/controller.extended_cond.opcode[1] ),
    .C(\heichips25_can_lehmann_fsm/_1145_ ),
    .A(\heichips25_can_lehmann_fsm/controller.extended_cond.opcode[2] ),
    .Y(\heichips25_can_lehmann_fsm/_1147_ ),
    .D(\heichips25_can_lehmann_fsm/_1146_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_1832_  (.A1(\heichips25_can_lehmann_fsm/net343 ),
    .A2(net4),
    .Y(\heichips25_can_lehmann_fsm/_1148_ ),
    .B1(\heichips25_can_lehmann_fsm/controller.extended_cond.opcode[1] ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_1833_  (.B1(\heichips25_can_lehmann_fsm/_1148_ ),
    .Y(\heichips25_can_lehmann_fsm/_1149_ ),
    .A1(\heichips25_can_lehmann_fsm/net343 ),
    .A2(\heichips25_can_lehmann_fsm/_0985_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_1834_  (.A1(\heichips25_can_lehmann_fsm/_1147_ ),
    .A2(\heichips25_can_lehmann_fsm/_1149_ ),
    .Y(\heichips25_can_lehmann_fsm/_1150_ ),
    .B1(\heichips25_can_lehmann_fsm/_1143_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_1835_  (.A1(\heichips25_can_lehmann_fsm/_1054_ ),
    .A2(\heichips25_can_lehmann_fsm/_1140_ ),
    .Y(\heichips25_can_lehmann_fsm/_1151_ ),
    .B1(\heichips25_can_lehmann_fsm/_1150_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_1836_  (.B1(\heichips25_can_lehmann_fsm/_1151_ ),
    .Y(\heichips25_can_lehmann_fsm/_1152_ ),
    .A1(\heichips25_can_lehmann_fsm/_1074_ ),
    .A2(\heichips25_can_lehmann_fsm/_1144_ ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_1837_  (.Y(\heichips25_can_lehmann_fsm/_1153_ ),
    .A(\heichips25_can_lehmann_fsm/net348 ),
    .B(\heichips25_can_lehmann_fsm/_0996_ ));
 sg13g2_xnor2_1 \heichips25_can_lehmann_fsm/_1838_  (.Y(\heichips25_can_lehmann_fsm/_1154_ ),
    .A(\heichips25_can_lehmann_fsm/controller.extended_state[1] ),
    .B(\heichips25_can_lehmann_fsm/net352 ));
 sg13g2_nand2b_1 \heichips25_can_lehmann_fsm/_1839_  (.Y(\heichips25_can_lehmann_fsm/_1155_ ),
    .B(\heichips25_can_lehmann_fsm/net348 ),
    .A_N(\heichips25_can_lehmann_fsm/controller.extended_state[2] ));
 sg13g2_xnor2_1 \heichips25_can_lehmann_fsm/_1840_  (.Y(\heichips25_can_lehmann_fsm/_1156_ ),
    .A(\heichips25_can_lehmann_fsm/controller.extended_state[0] ),
    .B(\heichips25_can_lehmann_fsm/net354 ));
 sg13g2_nand3_1 \heichips25_can_lehmann_fsm/_1841_  (.B(\heichips25_can_lehmann_fsm/_1155_ ),
    .C(\heichips25_can_lehmann_fsm/_1156_ ),
    .A(\heichips25_can_lehmann_fsm/_1154_ ),
    .Y(\heichips25_can_lehmann_fsm/_1157_ ));
 sg13g2_a21o_1 \heichips25_can_lehmann_fsm/_1842_  (.A2(\heichips25_can_lehmann_fsm/_1153_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.extended_state[2] ),
    .B1(\heichips25_can_lehmann_fsm/_1157_ ),
    .X(\heichips25_can_lehmann_fsm/_1158_ ));
 sg13g2_a21o_1 \heichips25_can_lehmann_fsm/_1843_  (.A2(\heichips25_can_lehmann_fsm/_1141_ ),
    .A1(\heichips25_can_lehmann_fsm/_1108_ ),
    .B1(\heichips25_can_lehmann_fsm/_1157_ ),
    .X(\heichips25_can_lehmann_fsm/_1159_ ));
 sg13g2_a21o_1 \heichips25_can_lehmann_fsm/_1844_  (.A2(\heichips25_can_lehmann_fsm/_1141_ ),
    .A1(\heichips25_can_lehmann_fsm/_1108_ ),
    .B1(\heichips25_can_lehmann_fsm/_1158_ ),
    .X(\heichips25_can_lehmann_fsm/_1160_ ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_1845_  (.B2(\heichips25_can_lehmann_fsm/controller.extended_state[2] ),
    .C1(\heichips25_can_lehmann_fsm/_1159_ ),
    .B1(\heichips25_can_lehmann_fsm/_1153_ ),
    .A1(\heichips25_can_lehmann_fsm/_1142_ ),
    .Y(\heichips25_can_lehmann_fsm/_1161_ ),
    .A2(\heichips25_can_lehmann_fsm/_1152_ ));
 sg13g2_a21o_1 \heichips25_can_lehmann_fsm/_1846_  (.A2(\heichips25_can_lehmann_fsm/_1152_ ),
    .A1(\heichips25_can_lehmann_fsm/_1142_ ),
    .B1(\heichips25_can_lehmann_fsm/_1160_ ),
    .X(\heichips25_can_lehmann_fsm/_1162_ ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_1847_  (.A(\heichips25_can_lehmann_fsm/_1139_ ),
    .B(\heichips25_can_lehmann_fsm/_1161_ ),
    .Y(\heichips25_can_lehmann_fsm/_1163_ ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1848_  (.Y(\heichips25_can_lehmann_fsm/_1164_ ),
    .A(\heichips25_can_lehmann_fsm/_1163_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_1849_  (.B1(\heichips25_can_lehmann_fsm/_1090_ ),
    .Y(\heichips25_can_lehmann_fsm/_1165_ ),
    .A1(\heichips25_can_lehmann_fsm/_1096_ ),
    .A2(\heichips25_can_lehmann_fsm/_1164_ ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_1850_  (.A(\heichips25_can_lehmann_fsm/_1139_ ),
    .B(\heichips25_can_lehmann_fsm/_1162_ ),
    .Y(\heichips25_can_lehmann_fsm/_1166_ ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1851_  (.Y(\heichips25_can_lehmann_fsm/_1167_ ),
    .B1(\heichips25_can_lehmann_fsm/net311 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[176] ),
    .A2(\heichips25_can_lehmann_fsm/net318 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[152] ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1852_  (.Y(\heichips25_can_lehmann_fsm/_1168_ ),
    .B1(\heichips25_can_lehmann_fsm/net297 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[56] ),
    .A2(\heichips25_can_lehmann_fsm/net307 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[104] ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1853_  (.Y(\heichips25_can_lehmann_fsm/_1169_ ),
    .B1(\heichips25_can_lehmann_fsm/net295 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[128] ),
    .A2(\heichips25_can_lehmann_fsm/net332 ),
    .A1(\heichips25_can_lehmann_fsm/controller.extended_jump_target[0] ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_1854_  (.A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[80] ),
    .A2(\heichips25_can_lehmann_fsm/net314 ),
    .Y(\heichips25_can_lehmann_fsm/_1170_ ),
    .B1(\heichips25_can_lehmann_fsm/net302 ));
 sg13g2_nand4_1 \heichips25_can_lehmann_fsm/_1855_  (.B(\heichips25_can_lehmann_fsm/_1168_ ),
    .C(\heichips25_can_lehmann_fsm/_1169_ ),
    .A(\heichips25_can_lehmann_fsm/_1167_ ),
    .Y(\heichips25_can_lehmann_fsm/_1171_ ),
    .D(\heichips25_can_lehmann_fsm/_1170_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_1856_  (.B1(\heichips25_can_lehmann_fsm/_1171_ ),
    .Y(\heichips25_can_lehmann_fsm/_1172_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[32] ),
    .A2(\heichips25_can_lehmann_fsm/net335 ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_1857_  (.A(\heichips25_can_lehmann_fsm/net219 ),
    .B(\heichips25_can_lehmann_fsm/_1172_ ),
    .Y(\heichips25_can_lehmann_fsm/_1173_ ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_1858_  (.B2(\heichips25_can_lehmann_fsm/net1160 ),
    .C1(\heichips25_can_lehmann_fsm/_1173_ ),
    .B1(\heichips25_can_lehmann_fsm/_1166_ ),
    .A1(\heichips25_can_lehmann_fsm/_0984_ ),
    .Y(\heichips25_can_lehmann_fsm/_1174_ ),
    .A2(\heichips25_can_lehmann_fsm/_1163_ ));
 sg13g2_nor2b_1 \heichips25_can_lehmann_fsm/_1859_  (.A(net9),
    .B_N(\heichips25_can_lehmann_fsm/net471 ),
    .Y(\heichips25_can_lehmann_fsm/_1175_ ));
 sg13g2_nand2b_1 \heichips25_can_lehmann_fsm/_1860_  (.Y(\heichips25_can_lehmann_fsm/_1176_ ),
    .B(\heichips25_can_lehmann_fsm/net471 ),
    .A_N(net9));
 sg13g2_mux2_1 \heichips25_can_lehmann_fsm/_1861_  (.A0(\heichips25_can_lehmann_fsm/_1174_ ),
    .A1(\heichips25_can_lehmann_fsm/_0984_ ),
    .S(\heichips25_can_lehmann_fsm/_1165_ ),
    .X(\heichips25_can_lehmann_fsm/_1177_ ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_1862_  (.A(\heichips25_can_lehmann_fsm/_1176_ ),
    .B(\heichips25_can_lehmann_fsm/_1177_ ),
    .Y(\heichips25_can_lehmann_fsm/_0000_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_1863_  (.A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[153] ),
    .A2(\heichips25_can_lehmann_fsm/net318 ),
    .Y(\heichips25_can_lehmann_fsm/_1178_ ),
    .B1(\heichips25_can_lehmann_fsm/net302 ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1864_  (.Y(\heichips25_can_lehmann_fsm/_1179_ ),
    .B1(\heichips25_can_lehmann_fsm/net332 ),
    .B2(\heichips25_can_lehmann_fsm/controller.extended_jump_target[1] ),
    .A2(\heichips25_can_lehmann_fsm/net307 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[105] ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1865_  (.Y(\heichips25_can_lehmann_fsm/_1180_ ),
    .B1(\heichips25_can_lehmann_fsm/net295 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[129] ),
    .A2(\heichips25_can_lehmann_fsm/net311 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[177] ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1866_  (.Y(\heichips25_can_lehmann_fsm/_1181_ ),
    .B1(\heichips25_can_lehmann_fsm/net297 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[57] ),
    .A2(\heichips25_can_lehmann_fsm/net314 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[81] ));
 sg13g2_nand4_1 \heichips25_can_lehmann_fsm/_1867_  (.B(\heichips25_can_lehmann_fsm/_1179_ ),
    .C(\heichips25_can_lehmann_fsm/_1180_ ),
    .A(\heichips25_can_lehmann_fsm/_1178_ ),
    .Y(\heichips25_can_lehmann_fsm/_1182_ ),
    .D(\heichips25_can_lehmann_fsm/_1181_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_1868_  (.B1(\heichips25_can_lehmann_fsm/_1182_ ),
    .Y(\heichips25_can_lehmann_fsm/_1183_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[33] ),
    .A2(\heichips25_can_lehmann_fsm/net335 ));
 sg13g2_nand3_1 \heichips25_can_lehmann_fsm/_1869_  (.B(\heichips25_can_lehmann_fsm/_0999_ ),
    .C(\heichips25_can_lehmann_fsm/_1163_ ),
    .A(\heichips25_can_lehmann_fsm/_0996_ ),
    .Y(\heichips25_can_lehmann_fsm/_1184_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_1870_  (.B1(\heichips25_can_lehmann_fsm/_1184_ ),
    .Y(\heichips25_can_lehmann_fsm/_1185_ ),
    .A1(\heichips25_can_lehmann_fsm/net219 ),
    .A2(\heichips25_can_lehmann_fsm/_1183_ ));
 sg13g2_a21o_1 \heichips25_can_lehmann_fsm/_1871_  (.A2(\heichips25_can_lehmann_fsm/_1166_ ),
    .A1(\heichips25_can_lehmann_fsm/net1172 ),
    .B1(\heichips25_can_lehmann_fsm/_1185_ ),
    .X(\heichips25_can_lehmann_fsm/_1186_ ));
 sg13g2_nand2b_1 \heichips25_can_lehmann_fsm/_1872_  (.Y(\heichips25_can_lehmann_fsm/_1187_ ),
    .B(\heichips25_can_lehmann_fsm/_1165_ ),
    .A_N(\heichips25_can_lehmann_fsm/net352 ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_1873_  (.B1(\heichips25_can_lehmann_fsm/_1187_ ),
    .Y(\heichips25_can_lehmann_fsm/_1188_ ),
    .A1(\heichips25_can_lehmann_fsm/_1165_ ),
    .A2(\heichips25_can_lehmann_fsm/_1186_ ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_1874_  (.A(\heichips25_can_lehmann_fsm/_1176_ ),
    .B(\heichips25_can_lehmann_fsm/_1188_ ),
    .Y(\heichips25_can_lehmann_fsm/_0001_ ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1875_  (.Y(\heichips25_can_lehmann_fsm/_1189_ ),
    .B1(\heichips25_can_lehmann_fsm/net307 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[106] ),
    .A2(\heichips25_can_lehmann_fsm/net311 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[178] ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1876_  (.Y(\heichips25_can_lehmann_fsm/_1190_ ),
    .B1(\heichips25_can_lehmann_fsm/net314 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[82] ),
    .A2(\heichips25_can_lehmann_fsm/net318 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[154] ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1877_  (.Y(\heichips25_can_lehmann_fsm/_1191_ ),
    .B1(\heichips25_can_lehmann_fsm/net295 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[130] ),
    .A2(\heichips25_can_lehmann_fsm/net332 ),
    .A1(\heichips25_can_lehmann_fsm/controller.extended_jump_target[2] ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_1878_  (.A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[58] ),
    .A2(\heichips25_can_lehmann_fsm/net297 ),
    .Y(\heichips25_can_lehmann_fsm/_1192_ ),
    .B1(\heichips25_can_lehmann_fsm/net302 ));
 sg13g2_nand4_1 \heichips25_can_lehmann_fsm/_1879_  (.B(\heichips25_can_lehmann_fsm/_1190_ ),
    .C(\heichips25_can_lehmann_fsm/_1191_ ),
    .A(\heichips25_can_lehmann_fsm/_1189_ ),
    .Y(\heichips25_can_lehmann_fsm/_1193_ ),
    .D(\heichips25_can_lehmann_fsm/_1192_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_1880_  (.B1(\heichips25_can_lehmann_fsm/_1193_ ),
    .Y(\heichips25_can_lehmann_fsm/_1194_ ),
    .A1(\heichips25_can_lehmann_fsm/net1272 ),
    .A2(\heichips25_can_lehmann_fsm/net335 ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_1881_  (.A(\heichips25_can_lehmann_fsm/net219 ),
    .B(\heichips25_can_lehmann_fsm/_1194_ ),
    .Y(\heichips25_can_lehmann_fsm/_1195_ ));
 sg13g2_nand2b_1 \heichips25_can_lehmann_fsm/_1882_  (.Y(\heichips25_can_lehmann_fsm/_1196_ ),
    .B(\heichips25_can_lehmann_fsm/_1153_ ),
    .A_N(\heichips25_can_lehmann_fsm/net305 ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_1883_  (.B2(\heichips25_can_lehmann_fsm/_1163_ ),
    .C1(\heichips25_can_lehmann_fsm/_1195_ ),
    .B1(\heichips25_can_lehmann_fsm/_1196_ ),
    .A1(\heichips25_can_lehmann_fsm/net1164 ),
    .Y(\heichips25_can_lehmann_fsm/_1197_ ),
    .A2(\heichips25_can_lehmann_fsm/_1166_ ));
 sg13g2_mux2_1 \heichips25_can_lehmann_fsm/_1884_  (.A0(\heichips25_can_lehmann_fsm/_1197_ ),
    .A1(\heichips25_can_lehmann_fsm/net338 ),
    .S(\heichips25_can_lehmann_fsm/_1165_ ),
    .X(\heichips25_can_lehmann_fsm/_1198_ ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_1885_  (.A(\heichips25_can_lehmann_fsm/_1176_ ),
    .B(\heichips25_can_lehmann_fsm/_1198_ ),
    .Y(\heichips25_can_lehmann_fsm/_0002_ ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_1886_  (.Y(\heichips25_can_lehmann_fsm/_1199_ ),
    .A(\heichips25_can_lehmann_fsm/_0941_ ),
    .B(\heichips25_can_lehmann_fsm/net302 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_1887_  (.A1(\heichips25_can_lehmann_fsm/_0893_ ),
    .A2(\heichips25_can_lehmann_fsm/net348 ),
    .Y(\heichips25_can_lehmann_fsm/_1200_ ),
    .B1(\heichips25_can_lehmann_fsm/_0999_ ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1888_  (.Y(\heichips25_can_lehmann_fsm/_1201_ ),
    .B1(\heichips25_can_lehmann_fsm/net307 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[125] ),
    .A2(\heichips25_can_lehmann_fsm/net311 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[197] ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1889_  (.Y(\heichips25_can_lehmann_fsm/_1202_ ),
    .B1(\heichips25_can_lehmann_fsm/net297 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[77] ),
    .A2(\heichips25_can_lehmann_fsm/net314 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[101] ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_1890_  (.B2(\heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[21] ),
    .C1(\heichips25_can_lehmann_fsm/_1200_ ),
    .B1(\heichips25_can_lehmann_fsm/net332 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[173] ),
    .Y(\heichips25_can_lehmann_fsm/_1203_ ),
    .A2(\heichips25_can_lehmann_fsm/net318 ));
 sg13g2_nand3_1 \heichips25_can_lehmann_fsm/_1891_  (.B(\heichips25_can_lehmann_fsm/_1202_ ),
    .C(\heichips25_can_lehmann_fsm/_1203_ ),
    .A(\heichips25_can_lehmann_fsm/_1201_ ),
    .Y(\heichips25_can_lehmann_fsm/_1204_ ));
 sg13g2_nand3_1 \heichips25_can_lehmann_fsm/_1892_  (.B(\heichips25_can_lehmann_fsm/_1199_ ),
    .C(\heichips25_can_lehmann_fsm/_1204_ ),
    .A(\heichips25_can_lehmann_fsm/_1162_ ),
    .Y(\heichips25_can_lehmann_fsm/_1205_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_1893_  (.A1(\heichips25_can_lehmann_fsm/controller.extended_then_action[3] ),
    .A2(\heichips25_can_lehmann_fsm/_1161_ ),
    .Y(\heichips25_can_lehmann_fsm/_1206_ ),
    .B1(\heichips25_can_lehmann_fsm/_1139_ ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_1894_  (.Y(\heichips25_can_lehmann_fsm/_1207_ ),
    .A(\heichips25_can_lehmann_fsm/_0896_ ),
    .B(\heichips25_can_lehmann_fsm/net349 ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1895_  (.Y(\heichips25_can_lehmann_fsm/_1208_ ),
    .B1(\heichips25_can_lehmann_fsm/_1207_ ),
    .B2(\heichips25_can_lehmann_fsm/net337 ),
    .A2(\heichips25_can_lehmann_fsm/net333 ),
    .A1(\heichips25_can_lehmann_fsm/controller.extended_then_action[3] ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1896_  (.Y(\heichips25_can_lehmann_fsm/_1209_ ),
    .B1(\heichips25_can_lehmann_fsm/net307 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[119] ),
    .A2(\heichips25_can_lehmann_fsm/net311 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[191] ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1897_  (.Y(\heichips25_can_lehmann_fsm/_1210_ ),
    .B1(\heichips25_can_lehmann_fsm/net314 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[95] ),
    .A2(\heichips25_can_lehmann_fsm/net318 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[167] ));
 sg13g2_nand3_1 \heichips25_can_lehmann_fsm/_1898_  (.B(\heichips25_can_lehmann_fsm/_1209_ ),
    .C(\heichips25_can_lehmann_fsm/_1210_ ),
    .A(\heichips25_can_lehmann_fsm/_1208_ ),
    .Y(\heichips25_can_lehmann_fsm/_1211_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_1899_  (.A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[71] ),
    .A2(\heichips25_can_lehmann_fsm/net297 ),
    .Y(\heichips25_can_lehmann_fsm/_1212_ ),
    .B1(\heichips25_can_lehmann_fsm/_1211_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_1900_  (.A1(\heichips25_can_lehmann_fsm/_0946_ ),
    .A2(\heichips25_can_lehmann_fsm/net302 ),
    .Y(\heichips25_can_lehmann_fsm/_1213_ ),
    .B1(\heichips25_can_lehmann_fsm/_1212_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_1901_  (.B1(\heichips25_can_lehmann_fsm/_1090_ ),
    .Y(\heichips25_can_lehmann_fsm/_1214_ ),
    .A1(\heichips25_can_lehmann_fsm/net219 ),
    .A2(\heichips25_can_lehmann_fsm/_1213_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_1902_  (.A1(\heichips25_can_lehmann_fsm/_1205_ ),
    .A2(\heichips25_can_lehmann_fsm/_1206_ ),
    .Y(\heichips25_can_lehmann_fsm/_1215_ ),
    .B1(\heichips25_can_lehmann_fsm/_1214_ ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_1903_  (.Y(\heichips25_can_lehmann_fsm/_1216_ ),
    .A(\heichips25_can_lehmann_fsm/_0940_ ),
    .B(\heichips25_can_lehmann_fsm/net302 ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_1904_  (.Y(\heichips25_can_lehmann_fsm/_1217_ ),
    .A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[175] ),
    .B(\heichips25_can_lehmann_fsm/net318 ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1905_  (.Y(\heichips25_can_lehmann_fsm/_1218_ ),
    .B1(\heichips25_can_lehmann_fsm/net307 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[127] ),
    .A2(\heichips25_can_lehmann_fsm/net311 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[199] ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1906_  (.Y(\heichips25_can_lehmann_fsm/_1219_ ),
    .B1(\heichips25_can_lehmann_fsm/net332 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[23] ),
    .A2(\heichips25_can_lehmann_fsm/net314 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[103] ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_1907_  (.Y(\heichips25_can_lehmann_fsm/_1220_ ),
    .A(\heichips25_can_lehmann_fsm/_0892_ ),
    .B(\heichips25_can_lehmann_fsm/net349 ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1908_  (.Y(\heichips25_can_lehmann_fsm/_1221_ ),
    .B1(\heichips25_can_lehmann_fsm/_1220_ ),
    .B2(\heichips25_can_lehmann_fsm/net337 ),
    .A2(\heichips25_can_lehmann_fsm/net297 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[79] ));
 sg13g2_nand4_1 \heichips25_can_lehmann_fsm/_1909_  (.B(\heichips25_can_lehmann_fsm/_1218_ ),
    .C(\heichips25_can_lehmann_fsm/_1219_ ),
    .A(\heichips25_can_lehmann_fsm/_1217_ ),
    .Y(\heichips25_can_lehmann_fsm/_1222_ ),
    .D(\heichips25_can_lehmann_fsm/_1221_ ));
 sg13g2_nand3_1 \heichips25_can_lehmann_fsm/_1910_  (.B(\heichips25_can_lehmann_fsm/_1216_ ),
    .C(\heichips25_can_lehmann_fsm/_1222_ ),
    .A(\heichips25_can_lehmann_fsm/_1162_ ),
    .Y(\heichips25_can_lehmann_fsm/_1223_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_1911_  (.A1(\heichips25_can_lehmann_fsm/controller.extended_then_action[5] ),
    .A2(\heichips25_can_lehmann_fsm/_1161_ ),
    .Y(\heichips25_can_lehmann_fsm/_1224_ ),
    .B1(\heichips25_can_lehmann_fsm/_1139_ ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_1912_  (.Y(\heichips25_can_lehmann_fsm/_1225_ ),
    .A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[97] ),
    .B(\heichips25_can_lehmann_fsm/net315 ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_1913_  (.Y(\heichips25_can_lehmann_fsm/_1226_ ),
    .A(\heichips25_can_lehmann_fsm/_0895_ ),
    .B(\heichips25_can_lehmann_fsm/net349 ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1914_  (.Y(\heichips25_can_lehmann_fsm/_1227_ ),
    .B1(\heichips25_can_lehmann_fsm/_1226_ ),
    .B2(\heichips25_can_lehmann_fsm/net337 ),
    .A2(\heichips25_can_lehmann_fsm/net297 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[73] ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1915_  (.Y(\heichips25_can_lehmann_fsm/_1228_ ),
    .B1(\heichips25_can_lehmann_fsm/net333 ),
    .B2(\heichips25_can_lehmann_fsm/controller.extended_then_action[5] ),
    .A2(\heichips25_can_lehmann_fsm/net308 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[121] ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1916_  (.Y(\heichips25_can_lehmann_fsm/_1229_ ),
    .B1(\heichips25_can_lehmann_fsm/net311 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[193] ),
    .A2(\heichips25_can_lehmann_fsm/net318 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[169] ));
 sg13g2_nand4_1 \heichips25_can_lehmann_fsm/_1917_  (.B(\heichips25_can_lehmann_fsm/_1227_ ),
    .C(\heichips25_can_lehmann_fsm/_1228_ ),
    .A(\heichips25_can_lehmann_fsm/_1225_ ),
    .Y(\heichips25_can_lehmann_fsm/_1230_ ),
    .D(\heichips25_can_lehmann_fsm/_1229_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_1918_  (.B1(\heichips25_can_lehmann_fsm/_1230_ ),
    .Y(\heichips25_can_lehmann_fsm/_1231_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[49] ),
    .A2(\heichips25_can_lehmann_fsm/net335 ));
 sg13g2_inv_1 \heichips25_can_lehmann_fsm/_1919_  (.Y(\heichips25_can_lehmann_fsm/_1232_ ),
    .A(\heichips25_can_lehmann_fsm/_1231_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_1920_  (.B1(\heichips25_can_lehmann_fsm/_1090_ ),
    .Y(\heichips25_can_lehmann_fsm/_1233_ ),
    .A1(\heichips25_can_lehmann_fsm/net219 ),
    .A2(\heichips25_can_lehmann_fsm/_1232_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_1921_  (.A1(\heichips25_can_lehmann_fsm/_1223_ ),
    .A2(\heichips25_can_lehmann_fsm/_1224_ ),
    .Y(\heichips25_can_lehmann_fsm/_1234_ ),
    .B1(\heichips25_can_lehmann_fsm/_1233_ ));
 sg13g2_a21o_1 \heichips25_can_lehmann_fsm/_1922_  (.A2(\heichips25_can_lehmann_fsm/_1224_ ),
    .A1(\heichips25_can_lehmann_fsm/_1223_ ),
    .B1(\heichips25_can_lehmann_fsm/_1233_ ),
    .X(\heichips25_can_lehmann_fsm/_1235_ ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_1923_  (.Y(\heichips25_can_lehmann_fsm/_1236_ ),
    .A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[126] ),
    .B(\heichips25_can_lehmann_fsm/net307 ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1924_  (.Y(\heichips25_can_lehmann_fsm/_1237_ ),
    .B1(\heichips25_can_lehmann_fsm/net314 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[102] ),
    .A2(\heichips25_can_lehmann_fsm/net318 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[174] ));
 sg13g2_nand2b_1 \heichips25_can_lehmann_fsm/_1925_  (.Y(\heichips25_can_lehmann_fsm/_1238_ ),
    .B(\heichips25_can_lehmann_fsm/net349 ),
    .A_N(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[150] ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1926_  (.Y(\heichips25_can_lehmann_fsm/_0289_ ),
    .B1(\heichips25_can_lehmann_fsm/net337 ),
    .B2(\heichips25_can_lehmann_fsm/_1238_ ),
    .A2(\heichips25_can_lehmann_fsm/net311 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[198] ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1927_  (.Y(\heichips25_can_lehmann_fsm/_0290_ ),
    .B1(\heichips25_can_lehmann_fsm/net332 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[22] ),
    .A2(\heichips25_can_lehmann_fsm/net297 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[78] ));
 sg13g2_nand4_1 \heichips25_can_lehmann_fsm/_1928_  (.B(\heichips25_can_lehmann_fsm/_1237_ ),
    .C(\heichips25_can_lehmann_fsm/_0289_ ),
    .A(\heichips25_can_lehmann_fsm/_1236_ ),
    .Y(\heichips25_can_lehmann_fsm/_0291_ ),
    .D(\heichips25_can_lehmann_fsm/_0290_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_1929_  (.B1(\heichips25_can_lehmann_fsm/_0291_ ),
    .Y(\heichips25_can_lehmann_fsm/_0292_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[54] ),
    .A2(\heichips25_can_lehmann_fsm/net336 ));
 sg13g2_nand2b_1 \heichips25_can_lehmann_fsm/_1930_  (.Y(\heichips25_can_lehmann_fsm/_0293_ ),
    .B(\heichips25_can_lehmann_fsm/_1162_ ),
    .A_N(\heichips25_can_lehmann_fsm/_0292_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_1931_  (.A1(\heichips25_can_lehmann_fsm/controller.extended_then_action[4] ),
    .A2(\heichips25_can_lehmann_fsm/_1161_ ),
    .Y(\heichips25_can_lehmann_fsm/_0294_ ),
    .B1(\heichips25_can_lehmann_fsm/_1139_ ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_1932_  (.Y(\heichips25_can_lehmann_fsm/_0295_ ),
    .A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[72] ),
    .B(\heichips25_can_lehmann_fsm/net298 ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_1933_  (.B1(\heichips25_can_lehmann_fsm/net337 ),
    .Y(\heichips25_can_lehmann_fsm/_0296_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[144] ),
    .A2(\heichips25_can_lehmann_fsm/net338 ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1934_  (.Y(\heichips25_can_lehmann_fsm/_0297_ ),
    .B1(\heichips25_can_lehmann_fsm/net333 ),
    .B2(\heichips25_can_lehmann_fsm/controller.extended_then_action[4] ),
    .A2(\heichips25_can_lehmann_fsm/net315 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[96] ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1935_  (.Y(\heichips25_can_lehmann_fsm/_0298_ ),
    .B1(\heichips25_can_lehmann_fsm/net312 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[192] ),
    .A2(\heichips25_can_lehmann_fsm/net319 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[168] ));
 sg13g2_nand4_1 \heichips25_can_lehmann_fsm/_1936_  (.B(\heichips25_can_lehmann_fsm/_0296_ ),
    .C(\heichips25_can_lehmann_fsm/_0297_ ),
    .A(\heichips25_can_lehmann_fsm/_0295_ ),
    .Y(\heichips25_can_lehmann_fsm/_0299_ ),
    .D(\heichips25_can_lehmann_fsm/_0298_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_1937_  (.A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[120] ),
    .A2(\heichips25_can_lehmann_fsm/net308 ),
    .Y(\heichips25_can_lehmann_fsm/_0300_ ),
    .B1(\heichips25_can_lehmann_fsm/_0299_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_1938_  (.A1(\heichips25_can_lehmann_fsm/_0945_ ),
    .A2(\heichips25_can_lehmann_fsm/net302 ),
    .Y(\heichips25_can_lehmann_fsm/_0301_ ),
    .B1(\heichips25_can_lehmann_fsm/_0300_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_1939_  (.B1(\heichips25_can_lehmann_fsm/_1090_ ),
    .Y(\heichips25_can_lehmann_fsm/_0302_ ),
    .A1(\heichips25_can_lehmann_fsm/net219 ),
    .A2(\heichips25_can_lehmann_fsm/_0301_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_1940_  (.A1(\heichips25_can_lehmann_fsm/_0293_ ),
    .A2(\heichips25_can_lehmann_fsm/_0294_ ),
    .Y(\heichips25_can_lehmann_fsm/_0303_ ),
    .B1(\heichips25_can_lehmann_fsm/_0302_ ));
 sg13g2_a21o_1 \heichips25_can_lehmann_fsm/_1941_  (.A2(\heichips25_can_lehmann_fsm/_0294_ ),
    .A1(\heichips25_can_lehmann_fsm/_0293_ ),
    .B1(\heichips25_can_lehmann_fsm/_0302_ ),
    .X(\heichips25_can_lehmann_fsm/_0304_ ));
 sg13g2_nor3_1 \heichips25_can_lehmann_fsm/_1942_  (.A(\heichips25_can_lehmann_fsm/_1215_ ),
    .B(\heichips25_can_lehmann_fsm/_1235_ ),
    .C(\heichips25_can_lehmann_fsm/_0304_ ),
    .Y(\heichips25_can_lehmann_fsm/_0305_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_1943_  (.A1(\heichips25_can_lehmann_fsm/_1215_ ),
    .A2(\heichips25_can_lehmann_fsm/_0303_ ),
    .Y(\heichips25_can_lehmann_fsm/_0306_ ),
    .B1(\heichips25_can_lehmann_fsm/_1234_ ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_1944_  (.A(\heichips25_can_lehmann_fsm/_1235_ ),
    .B(\heichips25_can_lehmann_fsm/_0303_ ),
    .Y(\heichips25_can_lehmann_fsm/_0307_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_1945_  (.A1(\heichips25_can_lehmann_fsm/net1253 ),
    .A2(\heichips25_can_lehmann_fsm/net188 ),
    .Y(\heichips25_can_lehmann_fsm/_0308_ ),
    .B1(\heichips25_can_lehmann_fsm/net192 ));
 sg13g2_and3_1 \heichips25_can_lehmann_fsm/_1946_  (.X(\heichips25_can_lehmann_fsm/_0309_ ),
    .A(\heichips25_can_lehmann_fsm/_1215_ ),
    .B(\heichips25_can_lehmann_fsm/_1234_ ),
    .C(\heichips25_can_lehmann_fsm/_0303_ ));
 sg13g2_xor2_1 \heichips25_can_lehmann_fsm/_1947_  (.B(\heichips25_can_lehmann_fsm/_1061_ ),
    .A(\heichips25_can_lehmann_fsm/net1242 ),
    .X(\heichips25_can_lehmann_fsm/_0310_ ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1948_  (.Y(\heichips25_can_lehmann_fsm/_0311_ ),
    .B1(\heichips25_can_lehmann_fsm/net186 ),
    .B2(\heichips25_can_lehmann_fsm/_0310_ ),
    .A2(\heichips25_can_lehmann_fsm/net199 ),
    .A1(\heichips25_can_lehmann_fsm/net1262 ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_1949_  (.A(\heichips25_can_lehmann_fsm/_1215_ ),
    .B(\heichips25_can_lehmann_fsm/_1234_ ),
    .Y(\heichips25_can_lehmann_fsm/_0312_ ));
 sg13g2_nand2b_1 \heichips25_can_lehmann_fsm/_1950_  (.Y(\heichips25_can_lehmann_fsm/_0313_ ),
    .B(\heichips25_can_lehmann_fsm/_1235_ ),
    .A_N(\heichips25_can_lehmann_fsm/_1215_ ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_1951_  (.A(\heichips25_can_lehmann_fsm/net347 ),
    .B(\heichips25_can_lehmann_fsm/net182 ),
    .Y(\heichips25_can_lehmann_fsm/_0314_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_1952_  (.B1(\heichips25_can_lehmann_fsm/net322 ),
    .Y(\heichips25_can_lehmann_fsm/_0315_ ),
    .A1(\heichips25_can_lehmann_fsm/net1242 ),
    .A2(\heichips25_can_lehmann_fsm/net179 ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_1953_  (.B2(\heichips25_can_lehmann_fsm/net195 ),
    .C1(\heichips25_can_lehmann_fsm/_0315_ ),
    .B1(\heichips25_can_lehmann_fsm/_0314_ ),
    .A1(\heichips25_can_lehmann_fsm/_0308_ ),
    .Y(\heichips25_can_lehmann_fsm/_0003_ ),
    .A2(\heichips25_can_lehmann_fsm/_0311_ ));
 sg13g2_xor2_1 \heichips25_can_lehmann_fsm/_1954_  (.B(\heichips25_can_lehmann_fsm/_1062_ ),
    .A(\heichips25_can_lehmann_fsm/net1253 ),
    .X(\heichips25_can_lehmann_fsm/_0316_ ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_1955_  (.Y(\heichips25_can_lehmann_fsm/_0317_ ),
    .A(\heichips25_can_lehmann_fsm/net184 ),
    .B(\heichips25_can_lehmann_fsm/_0316_ ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_1956_  (.B2(\heichips25_can_lehmann_fsm/net1249 ),
    .C1(\heichips25_can_lehmann_fsm/net191 ),
    .B1(\heichips25_can_lehmann_fsm/net188 ),
    .A1(\heichips25_can_lehmann_fsm/net1242 ),
    .Y(\heichips25_can_lehmann_fsm/_0318_ ),
    .A2(\heichips25_can_lehmann_fsm/net197 ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_1957_  (.B1(\heichips25_can_lehmann_fsm/net321 ),
    .Y(\heichips25_can_lehmann_fsm/_0319_ ),
    .A1(\heichips25_can_lehmann_fsm/net1253 ),
    .A2(\heichips25_can_lehmann_fsm/net178 ));
 sg13g2_nor2b_1 \heichips25_can_lehmann_fsm/_1958_  (.A(\heichips25_can_lehmann_fsm/net346 ),
    .B_N(\heichips25_can_lehmann_fsm/_1215_ ),
    .Y(\heichips25_can_lehmann_fsm/_0320_ ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_1959_  (.B2(\heichips25_can_lehmann_fsm/net191 ),
    .C1(\heichips25_can_lehmann_fsm/_0319_ ),
    .B1(\heichips25_can_lehmann_fsm/_0320_ ),
    .A1(\heichips25_can_lehmann_fsm/_0317_ ),
    .Y(\heichips25_can_lehmann_fsm/_0004_ ),
    .A2(\heichips25_can_lehmann_fsm/_0318_ ));
 sg13g2_xnor2_1 \heichips25_can_lehmann_fsm/_1960_  (.Y(\heichips25_can_lehmann_fsm/_0321_ ),
    .A(\heichips25_can_lehmann_fsm/net1249 ),
    .B(\heichips25_can_lehmann_fsm/_1063_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_1961_  (.A1(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[12] ),
    .A2(\heichips25_can_lehmann_fsm/net188 ),
    .Y(\heichips25_can_lehmann_fsm/_0322_ ),
    .B1(\heichips25_can_lehmann_fsm/net192 ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1962_  (.Y(\heichips25_can_lehmann_fsm/_0323_ ),
    .B1(\heichips25_can_lehmann_fsm/net184 ),
    .B2(\heichips25_can_lehmann_fsm/_0321_ ),
    .A2(\heichips25_can_lehmann_fsm/net197 ),
    .A1(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[10] ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_1963_  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[3] ),
    .B(\heichips25_can_lehmann_fsm/net181 ),
    .Y(\heichips25_can_lehmann_fsm/_0324_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_1964_  (.B1(\heichips25_can_lehmann_fsm/net322 ),
    .Y(\heichips25_can_lehmann_fsm/_0325_ ),
    .A1(\heichips25_can_lehmann_fsm/net1249 ),
    .A2(\heichips25_can_lehmann_fsm/net178 ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_1965_  (.B2(\heichips25_can_lehmann_fsm/net192 ),
    .C1(\heichips25_can_lehmann_fsm/_0325_ ),
    .B1(\heichips25_can_lehmann_fsm/_0324_ ),
    .A1(\heichips25_can_lehmann_fsm/_0322_ ),
    .Y(\heichips25_can_lehmann_fsm/_0005_ ),
    .A2(\heichips25_can_lehmann_fsm/_0323_ ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_1966_  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[12] ),
    .B(\heichips25_can_lehmann_fsm/_1065_ ),
    .Y(\heichips25_can_lehmann_fsm/_0326_ ));
 sg13g2_xnor2_1 \heichips25_can_lehmann_fsm/_1967_  (.Y(\heichips25_can_lehmann_fsm/_0327_ ),
    .A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[12] ),
    .B(\heichips25_can_lehmann_fsm/_1065_ ));
 sg13g2_and2_1 \heichips25_can_lehmann_fsm/_1968_  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[13] ),
    .B(\heichips25_can_lehmann_fsm/_0304_ ),
    .X(\heichips25_can_lehmann_fsm/_0328_ ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_1969_  (.B2(\heichips25_can_lehmann_fsm/_0327_ ),
    .C1(\heichips25_can_lehmann_fsm/_0328_ ),
    .B1(\heichips25_can_lehmann_fsm/net184 ),
    .A1(\heichips25_can_lehmann_fsm/net1249 ),
    .Y(\heichips25_can_lehmann_fsm/_0329_ ),
    .A2(\heichips25_can_lehmann_fsm/net197 ));
 sg13g2_or2_1 \heichips25_can_lehmann_fsm/_1970_  (.X(\heichips25_can_lehmann_fsm/_0330_ ),
    .B(\heichips25_can_lehmann_fsm/_0329_ ),
    .A(\heichips25_can_lehmann_fsm/net192 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_1971_  (.A1(\heichips25_can_lehmann_fsm/net345 ),
    .A2(\heichips25_can_lehmann_fsm/net192 ),
    .Y(\heichips25_can_lehmann_fsm/_0331_ ),
    .B1(\heichips25_can_lehmann_fsm/net181 ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_1972_  (.B1(\heichips25_can_lehmann_fsm/net322 ),
    .Y(\heichips25_can_lehmann_fsm/_0332_ ),
    .A1(\heichips25_can_lehmann_fsm/net1260 ),
    .A2(\heichips25_can_lehmann_fsm/net178 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_1973_  (.A1(\heichips25_can_lehmann_fsm/_0330_ ),
    .A2(\heichips25_can_lehmann_fsm/_0331_ ),
    .Y(\heichips25_can_lehmann_fsm/_0006_ ),
    .B1(\heichips25_can_lehmann_fsm/_0332_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_1974_  (.A1(\heichips25_can_lehmann_fsm/net1248 ),
    .A2(\heichips25_can_lehmann_fsm/net190 ),
    .Y(\heichips25_can_lehmann_fsm/_0333_ ),
    .B1(\heichips25_can_lehmann_fsm/net196 ));
 sg13g2_nor3_1 \heichips25_can_lehmann_fsm/_1975_  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[13] ),
    .B(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[12] ),
    .C(\heichips25_can_lehmann_fsm/_1065_ ),
    .Y(\heichips25_can_lehmann_fsm/_0334_ ));
 sg13g2_xor2_1 \heichips25_can_lehmann_fsm/_1976_  (.B(\heichips25_can_lehmann_fsm/_0326_ ),
    .A(\heichips25_can_lehmann_fsm/net1257 ),
    .X(\heichips25_can_lehmann_fsm/_0335_ ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1977_  (.Y(\heichips25_can_lehmann_fsm/_0336_ ),
    .B1(\heichips25_can_lehmann_fsm/net187 ),
    .B2(\heichips25_can_lehmann_fsm/_0335_ ),
    .A2(\heichips25_can_lehmann_fsm/net199 ),
    .A1(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[12] ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_1978_  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[5] ),
    .B(\heichips25_can_lehmann_fsm/net183 ),
    .Y(\heichips25_can_lehmann_fsm/_0337_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_1979_  (.B1(\heichips25_can_lehmann_fsm/net323 ),
    .Y(\heichips25_can_lehmann_fsm/_0338_ ),
    .A1(\heichips25_can_lehmann_fsm/net1257 ),
    .A2(\heichips25_can_lehmann_fsm/net179 ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_1980_  (.B2(\heichips25_can_lehmann_fsm/net196 ),
    .C1(\heichips25_can_lehmann_fsm/_0338_ ),
    .B1(\heichips25_can_lehmann_fsm/_0337_ ),
    .A1(\heichips25_can_lehmann_fsm/_0333_ ),
    .Y(\heichips25_can_lehmann_fsm/_0007_ ),
    .A2(\heichips25_can_lehmann_fsm/_0336_ ));
 sg13g2_nor2b_1 \heichips25_can_lehmann_fsm/_1981_  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[14] ),
    .B_N(\heichips25_can_lehmann_fsm/_0334_ ),
    .Y(\heichips25_can_lehmann_fsm/_0339_ ));
 sg13g2_nor2b_1 \heichips25_can_lehmann_fsm/_1982_  (.A(\heichips25_can_lehmann_fsm/_0334_ ),
    .B_N(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[14] ),
    .Y(\heichips25_can_lehmann_fsm/_0340_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_1983_  (.B1(\heichips25_can_lehmann_fsm/net185 ),
    .Y(\heichips25_can_lehmann_fsm/_0341_ ),
    .A1(\heichips25_can_lehmann_fsm/_0339_ ),
    .A2(\heichips25_can_lehmann_fsm/_0340_ ));
 sg13g2_nor2b_1 \heichips25_can_lehmann_fsm/_1984_  (.A(\heichips25_can_lehmann_fsm/net344 ),
    .B_N(\heichips25_can_lehmann_fsm/net193 ),
    .Y(\heichips25_can_lehmann_fsm/_0342_ ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_1985_  (.B2(\heichips25_can_lehmann_fsm/net1234 ),
    .C1(\heichips25_can_lehmann_fsm/net194 ),
    .B1(\heichips25_can_lehmann_fsm/net189 ),
    .A1(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[13] ),
    .Y(\heichips25_can_lehmann_fsm/_0343_ ),
    .A2(\heichips25_can_lehmann_fsm/net197 ));
 sg13g2_a21o_1 \heichips25_can_lehmann_fsm/_1986_  (.A2(\heichips25_can_lehmann_fsm/_0343_ ),
    .A1(\heichips25_can_lehmann_fsm/_0341_ ),
    .B1(\heichips25_can_lehmann_fsm/_0342_ ),
    .X(\heichips25_can_lehmann_fsm/_0344_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_1987_  (.B1(\heichips25_can_lehmann_fsm/net323 ),
    .Y(\heichips25_can_lehmann_fsm/_0345_ ),
    .A1(\heichips25_can_lehmann_fsm/net1248 ),
    .A2(\heichips25_can_lehmann_fsm/net177 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_1988_  (.A1(\heichips25_can_lehmann_fsm/net177 ),
    .A2(\heichips25_can_lehmann_fsm/_0344_ ),
    .Y(\heichips25_can_lehmann_fsm/_0008_ ),
    .B1(\heichips25_can_lehmann_fsm/_0345_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_1989_  (.A1(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[16] ),
    .A2(\heichips25_can_lehmann_fsm/net189 ),
    .Y(\heichips25_can_lehmann_fsm/_0346_ ),
    .B1(\heichips25_can_lehmann_fsm/net194 ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_1990_  (.B1(\heichips25_can_lehmann_fsm/_1067_ ),
    .Y(\heichips25_can_lehmann_fsm/_0347_ ),
    .A1(\heichips25_can_lehmann_fsm/_0982_ ),
    .A2(\heichips25_can_lehmann_fsm/_0339_ ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_1991_  (.Y(\heichips25_can_lehmann_fsm/_0348_ ),
    .B1(\heichips25_can_lehmann_fsm/net185 ),
    .B2(\heichips25_can_lehmann_fsm/_0347_ ),
    .A2(\heichips25_can_lehmann_fsm/net198 ),
    .A1(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[14] ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_1992_  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[7] ),
    .B(\heichips25_can_lehmann_fsm/net181 ),
    .Y(\heichips25_can_lehmann_fsm/_0349_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_1993_  (.B1(\heichips25_can_lehmann_fsm/net321 ),
    .Y(\heichips25_can_lehmann_fsm/_0350_ ),
    .A1(\heichips25_can_lehmann_fsm/net1234 ),
    .A2(\heichips25_can_lehmann_fsm/net177 ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_1994_  (.B2(\heichips25_can_lehmann_fsm/net194 ),
    .C1(\heichips25_can_lehmann_fsm/_0350_ ),
    .B1(\heichips25_can_lehmann_fsm/_0349_ ),
    .A1(\heichips25_can_lehmann_fsm/_0346_ ),
    .Y(\heichips25_can_lehmann_fsm/_0009_ ),
    .A2(\heichips25_can_lehmann_fsm/_0348_ ));
 sg13g2_xnor2_1 \heichips25_can_lehmann_fsm/_1995_  (.Y(\heichips25_can_lehmann_fsm/_0351_ ),
    .A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[16] ),
    .B(\heichips25_can_lehmann_fsm/_1067_ ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_1996_  (.Y(\heichips25_can_lehmann_fsm/_0352_ ),
    .A(\heichips25_can_lehmann_fsm/net185 ),
    .B(\heichips25_can_lehmann_fsm/_0351_ ));
 sg13g2_nor2b_1 \heichips25_can_lehmann_fsm/_1997_  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[8] ),
    .B_N(\heichips25_can_lehmann_fsm/net196 ),
    .Y(\heichips25_can_lehmann_fsm/_0353_ ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_1998_  (.B2(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[17] ),
    .C1(\heichips25_can_lehmann_fsm/net193 ),
    .B1(\heichips25_can_lehmann_fsm/net189 ),
    .A1(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[15] ),
    .Y(\heichips25_can_lehmann_fsm/_0354_ ),
    .A2(\heichips25_can_lehmann_fsm/net198 ));
 sg13g2_a21o_1 \heichips25_can_lehmann_fsm/_1999_  (.A2(\heichips25_can_lehmann_fsm/_0354_ ),
    .A1(\heichips25_can_lehmann_fsm/_0352_ ),
    .B1(\heichips25_can_lehmann_fsm/_0353_ ),
    .X(\heichips25_can_lehmann_fsm/_0355_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2000_  (.B1(\heichips25_can_lehmann_fsm/net326 ),
    .Y(\heichips25_can_lehmann_fsm/_0356_ ),
    .A1(\heichips25_can_lehmann_fsm/net1251 ),
    .A2(\heichips25_can_lehmann_fsm/net180 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2001_  (.A1(\heichips25_can_lehmann_fsm/net180 ),
    .A2(\heichips25_can_lehmann_fsm/_0355_ ),
    .Y(\heichips25_can_lehmann_fsm/_0010_ ),
    .B1(\heichips25_can_lehmann_fsm/_0356_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2002_  (.A1(\heichips25_can_lehmann_fsm/net1240 ),
    .A2(\heichips25_can_lehmann_fsm/net188 ),
    .Y(\heichips25_can_lehmann_fsm/_0357_ ),
    .B1(\heichips25_can_lehmann_fsm/net191 ));
 sg13g2_xnor2_1 \heichips25_can_lehmann_fsm/_2003_  (.Y(\heichips25_can_lehmann_fsm/_0358_ ),
    .A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[17] ),
    .B(\heichips25_can_lehmann_fsm/_1068_ ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_2004_  (.Y(\heichips25_can_lehmann_fsm/_0359_ ),
    .B1(\heichips25_can_lehmann_fsm/net184 ),
    .B2(\heichips25_can_lehmann_fsm/_0358_ ),
    .A2(\heichips25_can_lehmann_fsm/net197 ),
    .A1(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[16] ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_2005_  (.A(\heichips25_can_lehmann_fsm/net1242 ),
    .B(\heichips25_can_lehmann_fsm/net181 ),
    .Y(\heichips25_can_lehmann_fsm/_0360_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2006_  (.B1(\heichips25_can_lehmann_fsm/net321 ),
    .Y(\heichips25_can_lehmann_fsm/_0361_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[17] ),
    .A2(\heichips25_can_lehmann_fsm/net178 ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_2007_  (.B2(\heichips25_can_lehmann_fsm/net191 ),
    .C1(\heichips25_can_lehmann_fsm/_0361_ ),
    .B1(\heichips25_can_lehmann_fsm/_0360_ ),
    .A1(\heichips25_can_lehmann_fsm/_0357_ ),
    .Y(\heichips25_can_lehmann_fsm/_0011_ ),
    .A2(\heichips25_can_lehmann_fsm/_0359_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2008_  (.B1(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[18] ),
    .Y(\heichips25_can_lehmann_fsm/_0362_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[17] ),
    .A2(\heichips25_can_lehmann_fsm/_1068_ ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_2009_  (.Y(\heichips25_can_lehmann_fsm/_0363_ ),
    .A(\heichips25_can_lehmann_fsm/_1070_ ),
    .B(\heichips25_can_lehmann_fsm/_0362_ ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_2010_  (.Y(\heichips25_can_lehmann_fsm/_0364_ ),
    .A(\heichips25_can_lehmann_fsm/net184 ),
    .B(\heichips25_can_lehmann_fsm/_0363_ ));
 sg13g2_nor2b_1 \heichips25_can_lehmann_fsm/_2011_  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[10] ),
    .B_N(\heichips25_can_lehmann_fsm/net191 ),
    .Y(\heichips25_can_lehmann_fsm/_0365_ ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_2012_  (.B2(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[19] ),
    .C1(\heichips25_can_lehmann_fsm/net191 ),
    .B1(\heichips25_can_lehmann_fsm/net188 ),
    .A1(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[17] ),
    .Y(\heichips25_can_lehmann_fsm/_0366_ ),
    .A2(\heichips25_can_lehmann_fsm/net197 ));
 sg13g2_a21o_1 \heichips25_can_lehmann_fsm/_2013_  (.A2(\heichips25_can_lehmann_fsm/_0366_ ),
    .A1(\heichips25_can_lehmann_fsm/_0364_ ),
    .B1(\heichips25_can_lehmann_fsm/_0365_ ),
    .X(\heichips25_can_lehmann_fsm/_0367_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2014_  (.B1(\heichips25_can_lehmann_fsm/net321 ),
    .Y(\heichips25_can_lehmann_fsm/_0368_ ),
    .A1(\heichips25_can_lehmann_fsm/net1240 ),
    .A2(\heichips25_can_lehmann_fsm/net178 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2015_  (.A1(\heichips25_can_lehmann_fsm/net178 ),
    .A2(\heichips25_can_lehmann_fsm/_0367_ ),
    .Y(\heichips25_can_lehmann_fsm/_0012_ ),
    .B1(\heichips25_can_lehmann_fsm/_0368_ ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_2016_  (.B2(\heichips25_can_lehmann_fsm/net1246 ),
    .C1(\heichips25_can_lehmann_fsm/net181 ),
    .B1(\heichips25_can_lehmann_fsm/net188 ),
    .A1(\heichips25_can_lehmann_fsm/net1240 ),
    .Y(\heichips25_can_lehmann_fsm/_0369_ ),
    .A2(\heichips25_can_lehmann_fsm/net197 ));
 sg13g2_xnor2_1 \heichips25_can_lehmann_fsm/_2017_  (.Y(\heichips25_can_lehmann_fsm/_0370_ ),
    .A(\heichips25_can_lehmann_fsm/net1259 ),
    .B(\heichips25_can_lehmann_fsm/_1070_ ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_2018_  (.Y(\heichips25_can_lehmann_fsm/_0371_ ),
    .B1(\heichips25_can_lehmann_fsm/net184 ),
    .B2(\heichips25_can_lehmann_fsm/_0370_ ),
    .A2(\heichips25_can_lehmann_fsm/net191 ),
    .A1(\heichips25_can_lehmann_fsm/net1249 ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2019_  (.B1(\heichips25_can_lehmann_fsm/net321 ),
    .Y(\heichips25_can_lehmann_fsm/_0372_ ),
    .A1(\heichips25_can_lehmann_fsm/net1259 ),
    .A2(\heichips25_can_lehmann_fsm/net178 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2020_  (.A1(\heichips25_can_lehmann_fsm/_0369_ ),
    .A2(\heichips25_can_lehmann_fsm/_0371_ ),
    .Y(\heichips25_can_lehmann_fsm/_0013_ ),
    .B1(\heichips25_can_lehmann_fsm/_0372_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2021_  (.B1(\heichips25_can_lehmann_fsm/net1246 ),
    .Y(\heichips25_can_lehmann_fsm/_0373_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[19] ),
    .A2(\heichips25_can_lehmann_fsm/_1070_ ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_2022_  (.Y(\heichips25_can_lehmann_fsm/_0374_ ),
    .A(\heichips25_can_lehmann_fsm/_1072_ ),
    .B(\heichips25_can_lehmann_fsm/_0373_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2023_  (.A1(\heichips25_can_lehmann_fsm/net1244 ),
    .A2(\heichips25_can_lehmann_fsm/net188 ),
    .Y(\heichips25_can_lehmann_fsm/_0375_ ),
    .B1(\heichips25_can_lehmann_fsm/net191 ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_2024_  (.Y(\heichips25_can_lehmann_fsm/_0376_ ),
    .B1(\heichips25_can_lehmann_fsm/net184 ),
    .B2(\heichips25_can_lehmann_fsm/_0374_ ),
    .A2(\heichips25_can_lehmann_fsm/net197 ),
    .A1(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[19] ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_2025_  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[12] ),
    .B(\heichips25_can_lehmann_fsm/net181 ),
    .Y(\heichips25_can_lehmann_fsm/_0377_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2026_  (.B1(\heichips25_can_lehmann_fsm/net321 ),
    .Y(\heichips25_can_lehmann_fsm/_0378_ ),
    .A1(\heichips25_can_lehmann_fsm/net1246 ),
    .A2(\heichips25_can_lehmann_fsm/net178 ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_2027_  (.B2(\heichips25_can_lehmann_fsm/net192 ),
    .C1(\heichips25_can_lehmann_fsm/_0378_ ),
    .B1(\heichips25_can_lehmann_fsm/_0377_ ),
    .A1(\heichips25_can_lehmann_fsm/_0375_ ),
    .Y(\heichips25_can_lehmann_fsm/_0014_ ),
    .A2(\heichips25_can_lehmann_fsm/_0376_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2028_  (.A1(\heichips25_can_lehmann_fsm/net1238 ),
    .A2(\heichips25_can_lehmann_fsm/net189 ),
    .Y(\heichips25_can_lehmann_fsm/_0379_ ),
    .B1(\heichips25_can_lehmann_fsm/net193 ));
 sg13g2_xnor2_1 \heichips25_can_lehmann_fsm/_2029_  (.Y(\heichips25_can_lehmann_fsm/_0380_ ),
    .A(\heichips25_can_lehmann_fsm/_0980_ ),
    .B(\heichips25_can_lehmann_fsm/_1071_ ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_2030_  (.Y(\heichips25_can_lehmann_fsm/_0381_ ),
    .B1(\heichips25_can_lehmann_fsm/net185 ),
    .B2(\heichips25_can_lehmann_fsm/_0380_ ),
    .A2(\heichips25_can_lehmann_fsm/net198 ),
    .A1(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[20] ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_2031_  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[13] ),
    .B(\heichips25_can_lehmann_fsm/_0312_ ),
    .Y(\heichips25_can_lehmann_fsm/_0382_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2032_  (.B1(\heichips25_can_lehmann_fsm/net324 ),
    .Y(\heichips25_can_lehmann_fsm/_0383_ ),
    .A1(\heichips25_can_lehmann_fsm/net1244 ),
    .A2(\heichips25_can_lehmann_fsm/net177 ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_2033_  (.B2(\heichips25_can_lehmann_fsm/net193 ),
    .C1(\heichips25_can_lehmann_fsm/_0383_ ),
    .B1(\heichips25_can_lehmann_fsm/_0382_ ),
    .A1(\heichips25_can_lehmann_fsm/_0379_ ),
    .Y(\heichips25_can_lehmann_fsm/_0015_ ),
    .A2(\heichips25_can_lehmann_fsm/_0381_ ));
 sg13g2_xnor2_1 \heichips25_can_lehmann_fsm/_2034_  (.Y(\heichips25_can_lehmann_fsm/_0384_ ),
    .A(\heichips25_can_lehmann_fsm/_0979_ ),
    .B(\heichips25_can_lehmann_fsm/_1073_ ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_2035_  (.Y(\heichips25_can_lehmann_fsm/_0385_ ),
    .A(\heichips25_can_lehmann_fsm/net185 ),
    .B(\heichips25_can_lehmann_fsm/_0384_ ));
 sg13g2_nor2b_1 \heichips25_can_lehmann_fsm/_2036_  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[14] ),
    .B_N(\heichips25_can_lehmann_fsm/net193 ),
    .Y(\heichips25_can_lehmann_fsm/_0386_ ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_2037_  (.B2(\heichips25_can_lehmann_fsm/net1227 ),
    .C1(\heichips25_can_lehmann_fsm/net193 ),
    .B1(\heichips25_can_lehmann_fsm/net189 ),
    .A1(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[21] ),
    .Y(\heichips25_can_lehmann_fsm/_0387_ ),
    .A2(\heichips25_can_lehmann_fsm/net198 ));
 sg13g2_a21o_1 \heichips25_can_lehmann_fsm/_2038_  (.A2(\heichips25_can_lehmann_fsm/_0387_ ),
    .A1(\heichips25_can_lehmann_fsm/_0385_ ),
    .B1(\heichips25_can_lehmann_fsm/_0386_ ),
    .X(\heichips25_can_lehmann_fsm/_0388_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2039_  (.B1(\heichips25_can_lehmann_fsm/net324 ),
    .Y(\heichips25_can_lehmann_fsm/_0389_ ),
    .A1(\heichips25_can_lehmann_fsm/net1238 ),
    .A2(\heichips25_can_lehmann_fsm/net177 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2040_  (.A1(\heichips25_can_lehmann_fsm/net177 ),
    .A2(\heichips25_can_lehmann_fsm/_0388_ ),
    .Y(\heichips25_can_lehmann_fsm/_0016_ ),
    .B1(\heichips25_can_lehmann_fsm/_0389_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2041_  (.A1(\heichips25_can_lehmann_fsm/_0979_ ),
    .A2(\heichips25_can_lehmann_fsm/_1073_ ),
    .Y(\heichips25_can_lehmann_fsm/_0390_ ),
    .B1(\heichips25_can_lehmann_fsm/_0978_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2042_  (.B1(\heichips25_can_lehmann_fsm/net185 ),
    .Y(\heichips25_can_lehmann_fsm/_0391_ ),
    .A1(\heichips25_can_lehmann_fsm/_1074_ ),
    .A2(\heichips25_can_lehmann_fsm/_0390_ ));
 sg13g2_and2_1 \heichips25_can_lehmann_fsm/_2043_  (.A(net11),
    .B(\heichips25_can_lehmann_fsm/_1215_ ),
    .X(\heichips25_can_lehmann_fsm/_0392_ ));
 sg13g2_and2_1 \heichips25_can_lehmann_fsm/_2044_  (.A(\heichips25_can_lehmann_fsm/_0982_ ),
    .B(\heichips25_can_lehmann_fsm/net193 ),
    .X(\heichips25_can_lehmann_fsm/_0393_ ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_2045_  (.B2(\heichips25_can_lehmann_fsm/_0392_ ),
    .C1(\heichips25_can_lehmann_fsm/net193 ),
    .B1(\heichips25_can_lehmann_fsm/net189 ),
    .A1(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[22] ),
    .Y(\heichips25_can_lehmann_fsm/_0394_ ),
    .A2(\heichips25_can_lehmann_fsm/net198 ));
 sg13g2_a21o_1 \heichips25_can_lehmann_fsm/_2046_  (.A2(\heichips25_can_lehmann_fsm/_0394_ ),
    .A1(\heichips25_can_lehmann_fsm/_0391_ ),
    .B1(\heichips25_can_lehmann_fsm/_0393_ ),
    .X(\heichips25_can_lehmann_fsm/_0395_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2047_  (.B1(\heichips25_can_lehmann_fsm/net324 ),
    .Y(\heichips25_can_lehmann_fsm/_0396_ ),
    .A1(\heichips25_can_lehmann_fsm/net1227 ),
    .A2(\heichips25_can_lehmann_fsm/net177 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2048_  (.A1(\heichips25_can_lehmann_fsm/net177 ),
    .A2(\heichips25_can_lehmann_fsm/_0395_ ),
    .Y(\heichips25_can_lehmann_fsm/_0017_ ),
    .B1(\heichips25_can_lehmann_fsm/_0396_ ));
 sg13g2_xor2_1 \heichips25_can_lehmann_fsm/_2049_  (.B(\heichips25_can_lehmann_fsm/_1060_ ),
    .A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[8] ),
    .X(\heichips25_can_lehmann_fsm/_0397_ ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_2050_  (.Y(\heichips25_can_lehmann_fsm/_0398_ ),
    .B1(\heichips25_can_lehmann_fsm/net186 ),
    .B2(\heichips25_can_lehmann_fsm/_0397_ ),
    .A2(\heichips25_can_lehmann_fsm/net190 ),
    .A1(\heichips25_can_lehmann_fsm/net1242 ));
 sg13g2_xnor2_1 \heichips25_can_lehmann_fsm/_2051_  (.Y(\heichips25_can_lehmann_fsm/_0399_ ),
    .A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[3] ),
    .B(\heichips25_can_lehmann_fsm/net346 ));
 sg13g2_xor2_1 \heichips25_can_lehmann_fsm/_2052_  (.B(\heichips25_can_lehmann_fsm/net344 ),
    .A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[7] ),
    .X(\heichips25_can_lehmann_fsm/_0400_ ));
 sg13g2_xnor2_1 \heichips25_can_lehmann_fsm/_2053_  (.Y(\heichips25_can_lehmann_fsm/_0401_ ),
    .A(\heichips25_can_lehmann_fsm/_0399_ ),
    .B(\heichips25_can_lehmann_fsm/_0400_ ));
 sg13g2_xnor2_1 \heichips25_can_lehmann_fsm/_2054_  (.Y(\heichips25_can_lehmann_fsm/_0402_ ),
    .A(\heichips25_can_lehmann_fsm/net347 ),
    .B(\heichips25_can_lehmann_fsm/net1255 ));
 sg13g2_xnor2_1 \heichips25_can_lehmann_fsm/_2055_  (.Y(\heichips25_can_lehmann_fsm/_0403_ ),
    .A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[5] ),
    .B(\heichips25_can_lehmann_fsm/net345 ));
 sg13g2_xnor2_1 \heichips25_can_lehmann_fsm/_2056_  (.Y(\heichips25_can_lehmann_fsm/_0404_ ),
    .A(\heichips25_can_lehmann_fsm/_0402_ ),
    .B(\heichips25_can_lehmann_fsm/_0403_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2057_  (.B1(\heichips25_can_lehmann_fsm/_0303_ ),
    .Y(\heichips25_can_lehmann_fsm/_0405_ ),
    .A1(\heichips25_can_lehmann_fsm/_0401_ ),
    .A2(\heichips25_can_lehmann_fsm/_0404_ ));
 sg13g2_a21o_1 \heichips25_can_lehmann_fsm/_2058_  (.A2(\heichips25_can_lehmann_fsm/_0404_ ),
    .A1(\heichips25_can_lehmann_fsm/_0401_ ),
    .B1(\heichips25_can_lehmann_fsm/_0405_ ),
    .X(\heichips25_can_lehmann_fsm/_0406_ ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_2059_  (.Y(\heichips25_can_lehmann_fsm/_0407_ ),
    .B1(\heichips25_can_lehmann_fsm/net196 ),
    .B2(\heichips25_can_lehmann_fsm/_0406_ ),
    .A2(\heichips25_can_lehmann_fsm/net200 ),
    .A1(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[7] ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_2060_  (.A(\heichips25_can_lehmann_fsm/net1255 ),
    .B(\heichips25_can_lehmann_fsm/net182 ),
    .Y(\heichips25_can_lehmann_fsm/_0408_ ));
 sg13g2_nand2b_1 \heichips25_can_lehmann_fsm/_2061_  (.Y(\heichips25_can_lehmann_fsm/_0409_ ),
    .B(\heichips25_can_lehmann_fsm/_0304_ ),
    .A_N(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[8] ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2062_  (.B1(\heichips25_can_lehmann_fsm/net322 ),
    .Y(\heichips25_can_lehmann_fsm/_0410_ ),
    .A1(\heichips25_can_lehmann_fsm/net179 ),
    .A2(\heichips25_can_lehmann_fsm/_0409_ ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_2063_  (.B2(\heichips25_can_lehmann_fsm/net195 ),
    .C1(\heichips25_can_lehmann_fsm/_0410_ ),
    .B1(\heichips25_can_lehmann_fsm/_0408_ ),
    .A1(\heichips25_can_lehmann_fsm/_0398_ ),
    .Y(\heichips25_can_lehmann_fsm/_0018_ ),
    .A2(\heichips25_can_lehmann_fsm/_0407_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2064_  (.A1(\heichips25_can_lehmann_fsm/_1215_ ),
    .A2(\heichips25_can_lehmann_fsm/_0303_ ),
    .Y(\heichips25_can_lehmann_fsm/_0411_ ),
    .B1(\heichips25_can_lehmann_fsm/_0972_ ));
 sg13g2_nand2b_1 \heichips25_can_lehmann_fsm/_2065_  (.Y(\heichips25_can_lehmann_fsm/_0412_ ),
    .B(\heichips25_can_lehmann_fsm/_0411_ ),
    .A_N(\heichips25_can_lehmann_fsm/net189 ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_2066_  (.B2(\heichips25_can_lehmann_fsm/_0977_ ),
    .C1(\heichips25_can_lehmann_fsm/net181 ),
    .B1(\heichips25_can_lehmann_fsm/net184 ),
    .A1(\heichips25_can_lehmann_fsm/net347 ),
    .Y(\heichips25_can_lehmann_fsm/_0413_ ),
    .A2(\heichips25_can_lehmann_fsm/net188 ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_2067_  (.B2(\heichips25_can_lehmann_fsm/_0413_ ),
    .C1(\heichips25_can_lehmann_fsm/_1176_ ),
    .B1(\heichips25_can_lehmann_fsm/_0412_ ),
    .A1(\heichips25_can_lehmann_fsm/_0977_ ),
    .Y(\heichips25_can_lehmann_fsm/_0019_ ),
    .A2(\heichips25_can_lehmann_fsm/net181 ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_2068_  (.Y(\heichips25_can_lehmann_fsm/_0414_ ),
    .B1(\heichips25_can_lehmann_fsm/net186 ),
    .B2(\heichips25_can_lehmann_fsm/_0402_ ),
    .A2(\heichips25_can_lehmann_fsm/net195 ),
    .A1(net12));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_2069_  (.B2(\heichips25_can_lehmann_fsm/net346 ),
    .C1(\heichips25_can_lehmann_fsm/net182 ),
    .B1(\heichips25_can_lehmann_fsm/net190 ),
    .A1(\heichips25_can_lehmann_fsm/net1255 ),
    .Y(\heichips25_can_lehmann_fsm/_0415_ ),
    .A2(\heichips25_can_lehmann_fsm/net199 ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2070_  (.B1(\heichips25_can_lehmann_fsm/net322 ),
    .Y(\heichips25_can_lehmann_fsm/_0416_ ),
    .A1(\heichips25_can_lehmann_fsm/net347 ),
    .A2(\heichips25_can_lehmann_fsm/net179 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2071_  (.A1(\heichips25_can_lehmann_fsm/_0414_ ),
    .A2(\heichips25_can_lehmann_fsm/_0415_ ),
    .Y(\heichips25_can_lehmann_fsm/_0020_ ),
    .B1(\heichips25_can_lehmann_fsm/_0416_ ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_2072_  (.B2(\heichips25_can_lehmann_fsm/net1266 ),
    .C1(\heichips25_can_lehmann_fsm/net182 ),
    .B1(\heichips25_can_lehmann_fsm/net190 ),
    .A1(\heichips25_can_lehmann_fsm/net347 ),
    .Y(\heichips25_can_lehmann_fsm/_0417_ ),
    .A2(\heichips25_can_lehmann_fsm/net199 ));
 sg13g2_nor3_1 \heichips25_can_lehmann_fsm/_2073_  (.A(\heichips25_can_lehmann_fsm/net346 ),
    .B(\heichips25_can_lehmann_fsm/net347 ),
    .C(\heichips25_can_lehmann_fsm/net1274 ),
    .Y(\heichips25_can_lehmann_fsm/_0418_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2074_  (.B1(\heichips25_can_lehmann_fsm/net346 ),
    .Y(\heichips25_can_lehmann_fsm/_0419_ ),
    .A1(\heichips25_can_lehmann_fsm/net1269 ),
    .A2(\heichips25_can_lehmann_fsm/net1274 ));
 sg13g2_nand2b_1 \heichips25_can_lehmann_fsm/_2075_  (.Y(\heichips25_can_lehmann_fsm/_0420_ ),
    .B(\heichips25_can_lehmann_fsm/_0419_ ),
    .A_N(\heichips25_can_lehmann_fsm/_0418_ ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_2076_  (.Y(\heichips25_can_lehmann_fsm/_0421_ ),
    .B1(\heichips25_can_lehmann_fsm/net186 ),
    .B2(\heichips25_can_lehmann_fsm/_0420_ ),
    .A2(\heichips25_can_lehmann_fsm/net195 ),
    .A1(net13));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2077_  (.B1(\heichips25_can_lehmann_fsm/net322 ),
    .Y(\heichips25_can_lehmann_fsm/_0422_ ),
    .A1(\heichips25_can_lehmann_fsm/net346 ),
    .A2(\heichips25_can_lehmann_fsm/net179 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2078_  (.A1(\heichips25_can_lehmann_fsm/_0417_ ),
    .A2(\heichips25_can_lehmann_fsm/_0421_ ),
    .Y(\heichips25_can_lehmann_fsm/_0021_ ),
    .B1(\heichips25_can_lehmann_fsm/_0422_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2079_  (.B1(\heichips25_can_lehmann_fsm/_1056_ ),
    .Y(\heichips25_can_lehmann_fsm/_0423_ ),
    .A1(\heichips25_can_lehmann_fsm/_0976_ ),
    .A2(\heichips25_can_lehmann_fsm/_0418_ ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_2080_  (.B2(\heichips25_can_lehmann_fsm/_0423_ ),
    .C1(\heichips25_can_lehmann_fsm/net182 ),
    .B1(\heichips25_can_lehmann_fsm/net186 ),
    .A1(\heichips25_can_lehmann_fsm/net345 ),
    .Y(\heichips25_can_lehmann_fsm/_0424_ ),
    .A2(\heichips25_can_lehmann_fsm/net190 ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_2081_  (.Y(\heichips25_can_lehmann_fsm/_0425_ ),
    .B1(\heichips25_can_lehmann_fsm/net195 ),
    .B2(net14),
    .A2(\heichips25_can_lehmann_fsm/net199 ),
    .A1(\heichips25_can_lehmann_fsm/net1219 ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_2082_  (.B2(\heichips25_can_lehmann_fsm/_0425_ ),
    .C1(\heichips25_can_lehmann_fsm/_1176_ ),
    .B1(\heichips25_can_lehmann_fsm/_0424_ ),
    .A1(\heichips25_can_lehmann_fsm/_0976_ ),
    .Y(\heichips25_can_lehmann_fsm/_0022_ ),
    .A2(\heichips25_can_lehmann_fsm/net182 ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_2083_  (.B2(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[5] ),
    .C1(\heichips25_can_lehmann_fsm/net182 ),
    .B1(\heichips25_can_lehmann_fsm/net190 ),
    .A1(net15),
    .Y(\heichips25_can_lehmann_fsm/_0426_ ),
    .A2(\heichips25_can_lehmann_fsm/net195 ));
 sg13g2_xnor2_1 \heichips25_can_lehmann_fsm/_2084_  (.Y(\heichips25_can_lehmann_fsm/_0427_ ),
    .A(\heichips25_can_lehmann_fsm/net345 ),
    .B(\heichips25_can_lehmann_fsm/_1056_ ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_2085_  (.Y(\heichips25_can_lehmann_fsm/_0428_ ),
    .B1(\heichips25_can_lehmann_fsm/net186 ),
    .B2(\heichips25_can_lehmann_fsm/_0427_ ),
    .A2(\heichips25_can_lehmann_fsm/net199 ),
    .A1(\heichips25_can_lehmann_fsm/net1266 ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2086_  (.B1(\heichips25_can_lehmann_fsm/net322 ),
    .Y(\heichips25_can_lehmann_fsm/_0429_ ),
    .A1(\heichips25_can_lehmann_fsm/net345 ),
    .A2(\heichips25_can_lehmann_fsm/net179 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2087_  (.A1(\heichips25_can_lehmann_fsm/_0426_ ),
    .A2(\heichips25_can_lehmann_fsm/_0428_ ),
    .Y(\heichips25_can_lehmann_fsm/_0023_ ),
    .B1(\heichips25_can_lehmann_fsm/_0429_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2088_  (.B1(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[5] ),
    .Y(\heichips25_can_lehmann_fsm/_0430_ ),
    .A1(\heichips25_can_lehmann_fsm/net345 ),
    .A2(\heichips25_can_lehmann_fsm/_1056_ ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_2089_  (.Y(\heichips25_can_lehmann_fsm/_0431_ ),
    .A(\heichips25_can_lehmann_fsm/_1058_ ),
    .B(\heichips25_can_lehmann_fsm/_0430_ ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_2090_  (.Y(\heichips25_can_lehmann_fsm/_0432_ ),
    .A(\heichips25_can_lehmann_fsm/net186 ),
    .B(\heichips25_can_lehmann_fsm/_0431_ ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_2091_  (.Y(\heichips25_can_lehmann_fsm/_0433_ ),
    .B1(\heichips25_can_lehmann_fsm/net199 ),
    .B2(\heichips25_can_lehmann_fsm/net1264 ),
    .A2(\heichips25_can_lehmann_fsm/_0304_ ),
    .A1(\heichips25_can_lehmann_fsm/net344 ));
 sg13g2_a21o_1 \heichips25_can_lehmann_fsm/_2092_  (.A2(\heichips25_can_lehmann_fsm/_0433_ ),
    .A1(\heichips25_can_lehmann_fsm/_0432_ ),
    .B1(\heichips25_can_lehmann_fsm/net195 ),
    .X(\heichips25_can_lehmann_fsm/_0434_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2093_  (.A1(net16),
    .A2(\heichips25_can_lehmann_fsm/net195 ),
    .Y(\heichips25_can_lehmann_fsm/_0435_ ),
    .B1(\heichips25_can_lehmann_fsm/net182 ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2094_  (.B1(\heichips25_can_lehmann_fsm/net322 ),
    .Y(\heichips25_can_lehmann_fsm/_0436_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[5] ),
    .A2(\heichips25_can_lehmann_fsm/net179 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2095_  (.A1(\heichips25_can_lehmann_fsm/_0434_ ),
    .A2(\heichips25_can_lehmann_fsm/_0435_ ),
    .Y(\heichips25_can_lehmann_fsm/_0024_ ),
    .B1(\heichips25_can_lehmann_fsm/_0436_ ));
 sg13g2_xnor2_1 \heichips25_can_lehmann_fsm/_2096_  (.Y(\heichips25_can_lehmann_fsm/_0437_ ),
    .A(\heichips25_can_lehmann_fsm/net344 ),
    .B(\heichips25_can_lehmann_fsm/_1058_ ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_2097_  (.B2(\heichips25_can_lehmann_fsm/_0437_ ),
    .C1(\heichips25_can_lehmann_fsm/net183 ),
    .B1(\heichips25_can_lehmann_fsm/net186 ),
    .A1(\heichips25_can_lehmann_fsm/net1268 ),
    .Y(\heichips25_can_lehmann_fsm/_0438_ ),
    .A2(\heichips25_can_lehmann_fsm/_0307_ ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_2098_  (.Y(\heichips25_can_lehmann_fsm/_0439_ ),
    .B1(\heichips25_can_lehmann_fsm/net196 ),
    .B2(net17),
    .A2(\heichips25_can_lehmann_fsm/net199 ),
    .A1(\heichips25_can_lehmann_fsm/net1270 ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2099_  (.B1(\heichips25_can_lehmann_fsm/net323 ),
    .Y(\heichips25_can_lehmann_fsm/_0440_ ),
    .A1(\heichips25_can_lehmann_fsm/net344 ),
    .A2(\heichips25_can_lehmann_fsm/net179 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2100_  (.A1(\heichips25_can_lehmann_fsm/_0438_ ),
    .A2(\heichips25_can_lehmann_fsm/_0439_ ),
    .Y(\heichips25_can_lehmann_fsm/_0025_ ),
    .B1(\heichips25_can_lehmann_fsm/_0440_ ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_2101_  (.Y(\heichips25_can_lehmann_fsm/_0441_ ),
    .A(\heichips25_can_lehmann_fsm/net344 ),
    .B(\heichips25_can_lehmann_fsm/net200 ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2102_  (.B1(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[7] ),
    .Y(\heichips25_can_lehmann_fsm/_0442_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[6] ),
    .A2(\heichips25_can_lehmann_fsm/_1058_ ));
 sg13g2_nand2b_1 \heichips25_can_lehmann_fsm/_2103_  (.Y(\heichips25_can_lehmann_fsm/_0443_ ),
    .B(\heichips25_can_lehmann_fsm/_0442_ ),
    .A_N(\heichips25_can_lehmann_fsm/_1060_ ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_2104_  (.Y(\heichips25_can_lehmann_fsm/_0444_ ),
    .B1(\heichips25_can_lehmann_fsm/net187 ),
    .B2(\heichips25_can_lehmann_fsm/_0443_ ),
    .A2(\heichips25_can_lehmann_fsm/_0304_ ),
    .A1(\heichips25_can_lehmann_fsm/net1262 ));
 sg13g2_a21o_1 \heichips25_can_lehmann_fsm/_2105_  (.A2(\heichips25_can_lehmann_fsm/_0444_ ),
    .A1(\heichips25_can_lehmann_fsm/_0441_ ),
    .B1(\heichips25_can_lehmann_fsm/net196 ),
    .X(\heichips25_can_lehmann_fsm/_0445_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2106_  (.A1(net18),
    .A2(\heichips25_can_lehmann_fsm/net196 ),
    .Y(\heichips25_can_lehmann_fsm/_0446_ ),
    .B1(\heichips25_can_lehmann_fsm/net183 ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2107_  (.B1(\heichips25_can_lehmann_fsm/net323 ),
    .Y(\heichips25_can_lehmann_fsm/_0447_ ),
    .A1(\heichips25_can_lehmann_fsm/net1268 ),
    .A2(\heichips25_can_lehmann_fsm/net180 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2108_  (.A1(\heichips25_can_lehmann_fsm/_0445_ ),
    .A2(\heichips25_can_lehmann_fsm/_0446_ ),
    .Y(\heichips25_can_lehmann_fsm/_0026_ ),
    .B1(\heichips25_can_lehmann_fsm/_0447_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2109_  (.A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[195] ),
    .A2(\heichips25_can_lehmann_fsm/net312 ),
    .Y(\heichips25_can_lehmann_fsm/_0448_ ),
    .B1(\heichips25_can_lehmann_fsm/net303 ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_2110_  (.Y(\heichips25_can_lehmann_fsm/_0449_ ),
    .B1(\heichips25_can_lehmann_fsm/net298 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[75] ),
    .A2(\heichips25_can_lehmann_fsm/net308 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[123] ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_2111_  (.Y(\heichips25_can_lehmann_fsm/_0450_ ),
    .B1(\heichips25_can_lehmann_fsm/net295 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[147] ),
    .A2(\heichips25_can_lehmann_fsm/net315 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[99] ));
 sg13g2_nand3_1 \heichips25_can_lehmann_fsm/_2112_  (.B(\heichips25_can_lehmann_fsm/_0449_ ),
    .C(\heichips25_can_lehmann_fsm/_0450_ ),
    .A(\heichips25_can_lehmann_fsm/_0448_ ),
    .Y(\heichips25_can_lehmann_fsm/_0451_ ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_2113_  (.B2(\heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[19] ),
    .C1(\heichips25_can_lehmann_fsm/_0451_ ),
    .B1(\heichips25_can_lehmann_fsm/net333 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[171] ),
    .Y(\heichips25_can_lehmann_fsm/_0452_ ),
    .A2(\heichips25_can_lehmann_fsm/net319 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2114_  (.A1(\heichips25_can_lehmann_fsm/_0943_ ),
    .A2(\heichips25_can_lehmann_fsm/net303 ),
    .Y(\heichips25_can_lehmann_fsm/_0453_ ),
    .B1(\heichips25_can_lehmann_fsm/_0452_ ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_2115_  (.Y(\heichips25_can_lehmann_fsm/_0454_ ),
    .B1(\heichips25_can_lehmann_fsm/net331 ),
    .B2(\heichips25_can_lehmann_fsm/controller.extended_then_action[1] ),
    .A2(\heichips25_can_lehmann_fsm/net306 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[117] ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_2116_  (.Y(\heichips25_can_lehmann_fsm/_0455_ ),
    .B1(\heichips25_can_lehmann_fsm/net312 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[189] ),
    .A2(\heichips25_can_lehmann_fsm/net313 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[93] ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_2117_  (.Y(\heichips25_can_lehmann_fsm/_0456_ ),
    .B1(\heichips25_can_lehmann_fsm/net294 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[141] ),
    .A2(\heichips25_can_lehmann_fsm/net299 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[69] ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2118_  (.A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[165] ),
    .A2(\heichips25_can_lehmann_fsm/net317 ),
    .Y(\heichips25_can_lehmann_fsm/_0457_ ),
    .B1(\heichips25_can_lehmann_fsm/net301 ));
 sg13g2_nand4_1 \heichips25_can_lehmann_fsm/_2119_  (.B(\heichips25_can_lehmann_fsm/_0455_ ),
    .C(\heichips25_can_lehmann_fsm/_0456_ ),
    .A(\heichips25_can_lehmann_fsm/_0454_ ),
    .Y(\heichips25_can_lehmann_fsm/_0458_ ),
    .D(\heichips25_can_lehmann_fsm/_0457_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2120_  (.B1(\heichips25_can_lehmann_fsm/_0458_ ),
    .Y(\heichips25_can_lehmann_fsm/_0459_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[45] ),
    .A2(\heichips25_can_lehmann_fsm/net335 ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2121_  (.B1(\heichips25_can_lehmann_fsm/_1090_ ),
    .Y(\heichips25_can_lehmann_fsm/_0460_ ),
    .A1(\heichips25_can_lehmann_fsm/net219 ),
    .A2(\heichips25_can_lehmann_fsm/_0459_ ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_2122_  (.B2(\heichips25_can_lehmann_fsm/_1163_ ),
    .C1(\heichips25_can_lehmann_fsm/_0460_ ),
    .B1(\heichips25_can_lehmann_fsm/_0453_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.extended_then_action[1] ),
    .Y(\heichips25_can_lehmann_fsm/_0461_ ),
    .A2(\heichips25_can_lehmann_fsm/_1166_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2123_  (.A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[190] ),
    .A2(\heichips25_can_lehmann_fsm/net312 ),
    .Y(\heichips25_can_lehmann_fsm/_0462_ ),
    .B1(\heichips25_can_lehmann_fsm/net303 ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_2124_  (.Y(\heichips25_can_lehmann_fsm/_0463_ ),
    .B1(\heichips25_can_lehmann_fsm/net315 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[94] ),
    .A2(\heichips25_can_lehmann_fsm/net320 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[166] ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_2125_  (.Y(\heichips25_can_lehmann_fsm/_0464_ ),
    .B1(\heichips25_can_lehmann_fsm/net333 ),
    .B2(\heichips25_can_lehmann_fsm/controller.extended_then_action[2] ),
    .A2(\heichips25_can_lehmann_fsm/net299 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[70] ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_2126_  (.Y(\heichips25_can_lehmann_fsm/_0465_ ),
    .B1(\heichips25_can_lehmann_fsm/net295 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[142] ),
    .A2(\heichips25_can_lehmann_fsm/net306 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[118] ));
 sg13g2_nand4_1 \heichips25_can_lehmann_fsm/_2127_  (.B(\heichips25_can_lehmann_fsm/_0463_ ),
    .C(\heichips25_can_lehmann_fsm/_0464_ ),
    .A(\heichips25_can_lehmann_fsm/_0462_ ),
    .Y(\heichips25_can_lehmann_fsm/_0466_ ),
    .D(\heichips25_can_lehmann_fsm/_0465_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2128_  (.B1(\heichips25_can_lehmann_fsm/_0466_ ),
    .Y(\heichips25_can_lehmann_fsm/_0467_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[46] ),
    .A2(\heichips25_can_lehmann_fsm/net335 ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2129_  (.B1(\heichips25_can_lehmann_fsm/_1090_ ),
    .Y(\heichips25_can_lehmann_fsm/_0468_ ),
    .A1(\heichips25_can_lehmann_fsm/net219 ),
    .A2(\heichips25_can_lehmann_fsm/_0467_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2130_  (.B1(\heichips25_can_lehmann_fsm/net337 ),
    .Y(\heichips25_can_lehmann_fsm/_0469_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[148] ),
    .A2(\heichips25_can_lehmann_fsm/_0983_ ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_2131_  (.Y(\heichips25_can_lehmann_fsm/_0470_ ),
    .B1(\heichips25_can_lehmann_fsm/net332 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[20] ),
    .A2(\heichips25_can_lehmann_fsm/net319 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[172] ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_2132_  (.Y(\heichips25_can_lehmann_fsm/_0471_ ),
    .B1(\heichips25_can_lehmann_fsm/net307 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[124] ),
    .A2(\heichips25_can_lehmann_fsm/net315 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[100] ));
 sg13g2_nand3_1 \heichips25_can_lehmann_fsm/_2133_  (.B(\heichips25_can_lehmann_fsm/_0470_ ),
    .C(\heichips25_can_lehmann_fsm/_0471_ ),
    .A(\heichips25_can_lehmann_fsm/_0469_ ),
    .Y(\heichips25_can_lehmann_fsm/_0472_ ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_2134_  (.B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[76] ),
    .C1(\heichips25_can_lehmann_fsm/_0472_ ),
    .B1(\heichips25_can_lehmann_fsm/net298 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[196] ),
    .Y(\heichips25_can_lehmann_fsm/_0473_ ),
    .A2(\heichips25_can_lehmann_fsm/net312 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2135_  (.A1(\heichips25_can_lehmann_fsm/_0942_ ),
    .A2(\heichips25_can_lehmann_fsm/net303 ),
    .Y(\heichips25_can_lehmann_fsm/_0474_ ),
    .B1(\heichips25_can_lehmann_fsm/_0473_ ));
 sg13g2_mux2_1 \heichips25_can_lehmann_fsm/_2136_  (.A0(\heichips25_can_lehmann_fsm/controller.extended_then_action[2] ),
    .A1(\heichips25_can_lehmann_fsm/_0474_ ),
    .S(\heichips25_can_lehmann_fsm/_1162_ ),
    .X(\heichips25_can_lehmann_fsm/_0475_ ));
 sg13g2_a21o_1 \heichips25_can_lehmann_fsm/_2137_  (.A2(\heichips25_can_lehmann_fsm/_0475_ ),
    .A1(\heichips25_can_lehmann_fsm/_1138_ ),
    .B1(\heichips25_can_lehmann_fsm/_0468_ ),
    .X(\heichips25_can_lehmann_fsm/_0476_ ));
 sg13g2_nand2b_1 \heichips25_can_lehmann_fsm/_2138_  (.Y(\heichips25_can_lehmann_fsm/_0477_ ),
    .B(\heichips25_can_lehmann_fsm/net349 ),
    .A_N(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[146] ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_2139_  (.Y(\heichips25_can_lehmann_fsm/_0478_ ),
    .B1(\heichips25_can_lehmann_fsm/net308 ),
    .B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[122] ),
    .A2(\heichips25_can_lehmann_fsm/net319 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[170] ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_2140_  (.Y(\heichips25_can_lehmann_fsm/_0479_ ),
    .B1(\heichips25_can_lehmann_fsm/_0998_ ),
    .B2(\heichips25_can_lehmann_fsm/_0477_ ),
    .A2(\heichips25_can_lehmann_fsm/net315 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[98] ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2141_  (.B1(\heichips25_can_lehmann_fsm/_0479_ ),
    .Y(\heichips25_can_lehmann_fsm/_0480_ ),
    .A1(\heichips25_can_lehmann_fsm/_0868_ ),
    .A2(\heichips25_can_lehmann_fsm/_0995_ ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_2142_  (.B2(\heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[18] ),
    .C1(\heichips25_can_lehmann_fsm/_0480_ ),
    .B1(\heichips25_can_lehmann_fsm/net333 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[74] ),
    .Y(\heichips25_can_lehmann_fsm/_0481_ ),
    .A2(\heichips25_can_lehmann_fsm/net298 ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_2143_  (.Y(\heichips25_can_lehmann_fsm/_0482_ ),
    .B1(\heichips25_can_lehmann_fsm/_0478_ ),
    .B2(\heichips25_can_lehmann_fsm/_0481_ ),
    .A2(\heichips25_can_lehmann_fsm/net303 ),
    .A1(\heichips25_can_lehmann_fsm/_0944_ ));
 sg13g2_nand2b_1 \heichips25_can_lehmann_fsm/_2144_  (.Y(\heichips25_can_lehmann_fsm/_0483_ ),
    .B(\heichips25_can_lehmann_fsm/net348 ),
    .A_N(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[140] ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_2145_  (.Y(\heichips25_can_lehmann_fsm/_0484_ ),
    .B1(\heichips25_can_lehmann_fsm/net334 ),
    .B2(\heichips25_can_lehmann_fsm/controller.extended_then_action[0] ),
    .A2(\heichips25_can_lehmann_fsm/net299 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[68] ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_2146_  (.Y(\heichips25_can_lehmann_fsm/_0485_ ),
    .B1(\heichips25_can_lehmann_fsm/net337 ),
    .B2(\heichips25_can_lehmann_fsm/_0483_ ),
    .A2(\heichips25_can_lehmann_fsm/net316 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[92] ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2147_  (.B1(\heichips25_can_lehmann_fsm/_0485_ ),
    .Y(\heichips25_can_lehmann_fsm/_0486_ ),
    .A1(\heichips25_can_lehmann_fsm/_0884_ ),
    .A2(\heichips25_can_lehmann_fsm/_0991_ ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_2148_  (.B2(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[116] ),
    .C1(\heichips25_can_lehmann_fsm/_0486_ ),
    .B1(\heichips25_can_lehmann_fsm/net306 ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[188] ),
    .Y(\heichips25_can_lehmann_fsm/_0487_ ),
    .A2(\heichips25_can_lehmann_fsm/net312 ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_2149_  (.Y(\heichips25_can_lehmann_fsm/_0488_ ),
    .B1(\heichips25_can_lehmann_fsm/_0484_ ),
    .B2(\heichips25_can_lehmann_fsm/_0487_ ),
    .A2(\heichips25_can_lehmann_fsm/net301 ),
    .A1(\heichips25_can_lehmann_fsm/_0948_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2150_  (.B1(\heichips25_can_lehmann_fsm/_1090_ ),
    .Y(\heichips25_can_lehmann_fsm/_0489_ ),
    .A1(\heichips25_can_lehmann_fsm/_1138_ ),
    .A2(\heichips25_can_lehmann_fsm/_0488_ ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_2151_  (.Y(\heichips25_can_lehmann_fsm/_0490_ ),
    .A(\heichips25_can_lehmann_fsm/controller.extended_then_action[0] ),
    .B(\heichips25_can_lehmann_fsm/_1161_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2152_  (.A1(\heichips25_can_lehmann_fsm/_1162_ ),
    .A2(\heichips25_can_lehmann_fsm/_0482_ ),
    .Y(\heichips25_can_lehmann_fsm/_0491_ ),
    .B1(\heichips25_can_lehmann_fsm/_1139_ ));
 sg13g2_a21o_1 \heichips25_can_lehmann_fsm/_2153_  (.A2(\heichips25_can_lehmann_fsm/_0491_ ),
    .A1(\heichips25_can_lehmann_fsm/_0490_ ),
    .B1(\heichips25_can_lehmann_fsm/_0489_ ),
    .X(\heichips25_can_lehmann_fsm/_0492_ ));
 sg13g2_xnor2_1 \heichips25_can_lehmann_fsm/_2154_  (.Y(\heichips25_can_lehmann_fsm/_0493_ ),
    .A(\heichips25_can_lehmann_fsm/net205 ),
    .B(\heichips25_can_lehmann_fsm/_0492_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2155_  (.A1(\heichips25_can_lehmann_fsm/net205 ),
    .A2(\heichips25_can_lehmann_fsm/_0492_ ),
    .Y(\heichips25_can_lehmann_fsm/_0494_ ),
    .B1(\heichips25_can_lehmann_fsm/_0461_ ));
 sg13g2_a21o_1 \heichips25_can_lehmann_fsm/_2156_  (.A2(\heichips25_can_lehmann_fsm/_0492_ ),
    .A1(\heichips25_can_lehmann_fsm/net205 ),
    .B1(\heichips25_can_lehmann_fsm/_0461_ ),
    .X(\heichips25_can_lehmann_fsm/_0495_ ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_2157_  (.A(\heichips25_can_lehmann_fsm/_0461_ ),
    .B(\heichips25_can_lehmann_fsm/_0493_ ),
    .Y(\heichips25_can_lehmann_fsm/_0496_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2158_  (.A1(\heichips25_can_lehmann_fsm/_0461_ ),
    .A2(\heichips25_can_lehmann_fsm/_0493_ ),
    .Y(\heichips25_can_lehmann_fsm/_0497_ ),
    .B1(\heichips25_can_lehmann_fsm/_0494_ ));
 sg13g2_a21o_1 \heichips25_can_lehmann_fsm/_2159_  (.A2(\heichips25_can_lehmann_fsm/_0493_ ),
    .A1(\heichips25_can_lehmann_fsm/_0461_ ),
    .B1(\heichips25_can_lehmann_fsm/_0494_ ),
    .X(\heichips25_can_lehmann_fsm/_0498_ ));
 sg13g2_nor3_1 \heichips25_can_lehmann_fsm/_2160_  (.A(\heichips25_can_lehmann_fsm/_0461_ ),
    .B(\heichips25_can_lehmann_fsm/net205 ),
    .C(\heichips25_can_lehmann_fsm/_0492_ ),
    .Y(\heichips25_can_lehmann_fsm/_0499_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2161_  (.A1(net11),
    .A2(\heichips25_can_lehmann_fsm/_0499_ ),
    .Y(\heichips25_can_lehmann_fsm/_0500_ ),
    .B1(\heichips25_can_lehmann_fsm/_0497_ ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_2162_  (.Y(\heichips25_can_lehmann_fsm/_0501_ ),
    .B1(\heichips25_can_lehmann_fsm/net164 ),
    .B2(\heichips25_can_lehmann_fsm/_0975_ ),
    .A2(\heichips25_can_lehmann_fsm/net175 ),
    .A1(\heichips25_can_lehmann_fsm/net1204 ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_2163_  (.B2(\heichips25_can_lehmann_fsm/_0501_ ),
    .C1(\heichips25_can_lehmann_fsm/_1176_ ),
    .B1(\heichips25_can_lehmann_fsm/_0500_ ),
    .A1(\heichips25_can_lehmann_fsm/_0975_ ),
    .Y(\heichips25_can_lehmann_fsm/_0027_ ),
    .A2(\heichips25_can_lehmann_fsm/_0497_ ));
 sg13g2_xnor2_1 \heichips25_can_lehmann_fsm/_2164_  (.Y(\heichips25_can_lehmann_fsm/_0502_ ),
    .A(\heichips25_can_lehmann_fsm/net1233 ),
    .B(\heichips25_can_lehmann_fsm/net1226 ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_2165_  (.Y(\heichips25_can_lehmann_fsm/_0503_ ),
    .A(\heichips25_can_lehmann_fsm/net164 ),
    .B(\heichips25_can_lehmann_fsm/_0502_ ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_2166_  (.B2(net12),
    .C1(\heichips25_can_lehmann_fsm/_0497_ ),
    .B1(\heichips25_can_lehmann_fsm/_0499_ ),
    .A1(\heichips25_can_lehmann_fsm/net1093 ),
    .Y(\heichips25_can_lehmann_fsm/_0504_ ),
    .A2(\heichips25_can_lehmann_fsm/net175 ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2167_  (.B1(\heichips25_can_lehmann_fsm/net325 ),
    .Y(\heichips25_can_lehmann_fsm/_0505_ ),
    .A1(\heichips25_can_lehmann_fsm/net1233 ),
    .A2(\heichips25_can_lehmann_fsm/net160 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2168_  (.A1(\heichips25_can_lehmann_fsm/_0503_ ),
    .A2(\heichips25_can_lehmann_fsm/_0504_ ),
    .Y(\heichips25_can_lehmann_fsm/_0028_ ),
    .B1(\heichips25_can_lehmann_fsm/_0505_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2169_  (.B1(\heichips25_can_lehmann_fsm/net1215 ),
    .Y(\heichips25_can_lehmann_fsm/_0506_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[1] ),
    .A2(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[0] ));
 sg13g2_nand2b_1 \heichips25_can_lehmann_fsm/_2170_  (.Y(\heichips25_can_lehmann_fsm/_0507_ ),
    .B(\heichips25_can_lehmann_fsm/_0506_ ),
    .A_N(\heichips25_can_lehmann_fsm/_1097_ ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_2171_  (.Y(\heichips25_can_lehmann_fsm/_0508_ ),
    .A(\heichips25_can_lehmann_fsm/net164 ),
    .B(\heichips25_can_lehmann_fsm/_0507_ ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_2172_  (.B2(net13),
    .C1(\heichips25_can_lehmann_fsm/_0497_ ),
    .B1(\heichips25_can_lehmann_fsm/_0499_ ),
    .A1(\heichips25_can_lehmann_fsm/net1136 ),
    .Y(\heichips25_can_lehmann_fsm/_0509_ ),
    .A2(\heichips25_can_lehmann_fsm/net175 ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2173_  (.B1(\heichips25_can_lehmann_fsm/net325 ),
    .Y(\heichips25_can_lehmann_fsm/_0510_ ),
    .A1(\heichips25_can_lehmann_fsm/net1215 ),
    .A2(\heichips25_can_lehmann_fsm/net160 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2174_  (.A1(\heichips25_can_lehmann_fsm/_0508_ ),
    .A2(\heichips25_can_lehmann_fsm/_0509_ ),
    .Y(\heichips25_can_lehmann_fsm/_0029_ ),
    .B1(\heichips25_can_lehmann_fsm/_0510_ ));
 sg13g2_xor2_1 \heichips25_can_lehmann_fsm/_2175_  (.B(\heichips25_can_lehmann_fsm/_1097_ ),
    .A(\heichips25_can_lehmann_fsm/net1202 ),
    .X(\heichips25_can_lehmann_fsm/_0511_ ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_2176_  (.A(\heichips25_can_lehmann_fsm/_0970_ ),
    .B(\heichips25_can_lehmann_fsm/_0494_ ),
    .Y(\heichips25_can_lehmann_fsm/_0512_ ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_2177_  (.B2(\heichips25_can_lehmann_fsm/net164 ),
    .C1(\heichips25_can_lehmann_fsm/_0512_ ),
    .B1(\heichips25_can_lehmann_fsm/_0511_ ),
    .A1(net14),
    .Y(\heichips25_can_lehmann_fsm/_0513_ ),
    .A2(\heichips25_can_lehmann_fsm/_0499_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2178_  (.B1(\heichips25_can_lehmann_fsm/net325 ),
    .Y(\heichips25_can_lehmann_fsm/_0514_ ),
    .A1(\heichips25_can_lehmann_fsm/net1202 ),
    .A2(\heichips25_can_lehmann_fsm/net160 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2179_  (.A1(\heichips25_can_lehmann_fsm/net160 ),
    .A2(\heichips25_can_lehmann_fsm/_0513_ ),
    .Y(\heichips25_can_lehmann_fsm/_0030_ ),
    .B1(\heichips25_can_lehmann_fsm/_0514_ ));
 sg13g2_xnor2_1 \heichips25_can_lehmann_fsm/_2180_  (.Y(\heichips25_can_lehmann_fsm/_0515_ ),
    .A(\heichips25_can_lehmann_fsm/net1236 ),
    .B(\heichips25_can_lehmann_fsm/_1098_ ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_2181_  (.Y(\heichips25_can_lehmann_fsm/_0516_ ),
    .A(\heichips25_can_lehmann_fsm/net164 ),
    .B(\heichips25_can_lehmann_fsm/_0515_ ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_2182_  (.B2(net15),
    .C1(\heichips25_can_lehmann_fsm/_0497_ ),
    .B1(\heichips25_can_lehmann_fsm/_0499_ ),
    .A1(\heichips25_can_lehmann_fsm/net933 ),
    .Y(\heichips25_can_lehmann_fsm/_0517_ ),
    .A2(\heichips25_can_lehmann_fsm/net175 ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2183_  (.B1(\heichips25_can_lehmann_fsm/net325 ),
    .Y(\heichips25_can_lehmann_fsm/_0518_ ),
    .A1(\heichips25_can_lehmann_fsm/net1236 ),
    .A2(\heichips25_can_lehmann_fsm/net160 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2184_  (.A1(\heichips25_can_lehmann_fsm/_0516_ ),
    .A2(\heichips25_can_lehmann_fsm/_0517_ ),
    .Y(\heichips25_can_lehmann_fsm/_0031_ ),
    .B1(\heichips25_can_lehmann_fsm/_0518_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2185_  (.B1(\heichips25_can_lehmann_fsm/net1210 ),
    .Y(\heichips25_can_lehmann_fsm/_0519_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[4] ),
    .A2(\heichips25_can_lehmann_fsm/_1098_ ));
 sg13g2_nand2b_1 \heichips25_can_lehmann_fsm/_2186_  (.Y(\heichips25_can_lehmann_fsm/_0520_ ),
    .B(\heichips25_can_lehmann_fsm/_0519_ ),
    .A_N(\heichips25_can_lehmann_fsm/_1099_ ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_2187_  (.A(\heichips25_can_lehmann_fsm/_0969_ ),
    .B(\heichips25_can_lehmann_fsm/_0494_ ),
    .Y(\heichips25_can_lehmann_fsm/_0521_ ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_2188_  (.B2(\heichips25_can_lehmann_fsm/net164 ),
    .C1(\heichips25_can_lehmann_fsm/_0521_ ),
    .B1(\heichips25_can_lehmann_fsm/_0520_ ),
    .A1(net16),
    .Y(\heichips25_can_lehmann_fsm/_0522_ ),
    .A2(\heichips25_can_lehmann_fsm/_0499_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2189_  (.B1(\heichips25_can_lehmann_fsm/net325 ),
    .Y(\heichips25_can_lehmann_fsm/_0523_ ),
    .A1(\heichips25_can_lehmann_fsm/net1210 ),
    .A2(\heichips25_can_lehmann_fsm/net160 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2190_  (.A1(\heichips25_can_lehmann_fsm/net160 ),
    .A2(\heichips25_can_lehmann_fsm/_0522_ ),
    .Y(\heichips25_can_lehmann_fsm/_0032_ ),
    .B1(\heichips25_can_lehmann_fsm/_0523_ ));
 sg13g2_nor2b_1 \heichips25_can_lehmann_fsm/_2191_  (.A(\heichips25_can_lehmann_fsm/_1099_ ),
    .B_N(\heichips25_can_lehmann_fsm/net1192 ),
    .Y(\heichips25_can_lehmann_fsm/_0524_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2192_  (.B1(\heichips25_can_lehmann_fsm/net164 ),
    .Y(\heichips25_can_lehmann_fsm/_0525_ ),
    .A1(\heichips25_can_lehmann_fsm/_1100_ ),
    .A2(\heichips25_can_lehmann_fsm/_0524_ ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_2193_  (.B2(net17),
    .C1(\heichips25_can_lehmann_fsm/_0497_ ),
    .B1(\heichips25_can_lehmann_fsm/_0499_ ),
    .A1(\heichips25_can_lehmann_fsm/net1113 ),
    .Y(\heichips25_can_lehmann_fsm/_0526_ ),
    .A2(\heichips25_can_lehmann_fsm/net175 ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2194_  (.B1(\heichips25_can_lehmann_fsm/net325 ),
    .Y(\heichips25_can_lehmann_fsm/_0527_ ),
    .A1(\heichips25_can_lehmann_fsm/net1192 ),
    .A2(\heichips25_can_lehmann_fsm/net160 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2195_  (.A1(\heichips25_can_lehmann_fsm/_0525_ ),
    .A2(\heichips25_can_lehmann_fsm/_0526_ ),
    .Y(\heichips25_can_lehmann_fsm/_0033_ ),
    .B1(\heichips25_can_lehmann_fsm/_0527_ ));
 sg13g2_xnor2_1 \heichips25_can_lehmann_fsm/_2196_  (.Y(\heichips25_can_lehmann_fsm/_0528_ ),
    .A(\heichips25_can_lehmann_fsm/_0974_ ),
    .B(\heichips25_can_lehmann_fsm/_1100_ ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_2197_  (.Y(\heichips25_can_lehmann_fsm/_0529_ ),
    .A(\heichips25_can_lehmann_fsm/net164 ),
    .B(\heichips25_can_lehmann_fsm/_0528_ ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_2198_  (.B2(net18),
    .C1(\heichips25_can_lehmann_fsm/_0497_ ),
    .B1(\heichips25_can_lehmann_fsm/_0499_ ),
    .A1(\heichips25_can_lehmann_fsm/net1088 ),
    .Y(\heichips25_can_lehmann_fsm/_0530_ ),
    .A2(\heichips25_can_lehmann_fsm/net175 ));
 sg13g2_a221oi_1 \heichips25_can_lehmann_fsm/_2199_  (.B2(\heichips25_can_lehmann_fsm/_0530_ ),
    .C1(\heichips25_can_lehmann_fsm/_1176_ ),
    .B1(\heichips25_can_lehmann_fsm/_0529_ ),
    .A1(\heichips25_can_lehmann_fsm/_0974_ ),
    .Y(\heichips25_can_lehmann_fsm/_0034_ ),
    .A2(\heichips25_can_lehmann_fsm/_0497_ ));
 sg13g2_xnor2_1 \heichips25_can_lehmann_fsm/_2200_  (.Y(\heichips25_can_lehmann_fsm/_0531_ ),
    .A(\heichips25_can_lehmann_fsm/net1218 ),
    .B(\heichips25_can_lehmann_fsm/_1101_ ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_2201_  (.Y(\heichips25_can_lehmann_fsm/_0532_ ),
    .B1(\heichips25_can_lehmann_fsm/net165 ),
    .B2(\heichips25_can_lehmann_fsm/_0531_ ),
    .A2(\heichips25_can_lehmann_fsm/net175 ),
    .A1(\heichips25_can_lehmann_fsm/net974 ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2202_  (.B1(\heichips25_can_lehmann_fsm/net325 ),
    .Y(\heichips25_can_lehmann_fsm/_0533_ ),
    .A1(\heichips25_can_lehmann_fsm/net1218 ),
    .A2(\heichips25_can_lehmann_fsm/net163 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2203_  (.A1(\heichips25_can_lehmann_fsm/net163 ),
    .A2(\heichips25_can_lehmann_fsm/_0532_ ),
    .Y(\heichips25_can_lehmann_fsm/_0035_ ),
    .B1(\heichips25_can_lehmann_fsm/_0533_ ));
 sg13g2_xnor2_1 \heichips25_can_lehmann_fsm/_2204_  (.Y(\heichips25_can_lehmann_fsm/_0534_ ),
    .A(\heichips25_can_lehmann_fsm/net1180 ),
    .B(\heichips25_can_lehmann_fsm/_1102_ ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_2205_  (.Y(\heichips25_can_lehmann_fsm/_0535_ ),
    .B1(\heichips25_can_lehmann_fsm/net165 ),
    .B2(\heichips25_can_lehmann_fsm/_0534_ ),
    .A2(\heichips25_can_lehmann_fsm/net175 ),
    .A1(\heichips25_can_lehmann_fsm/net851 ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2206_  (.B1(\heichips25_can_lehmann_fsm/net325 ),
    .Y(\heichips25_can_lehmann_fsm/_0536_ ),
    .A1(\heichips25_can_lehmann_fsm/net1180 ),
    .A2(\heichips25_can_lehmann_fsm/net161 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2207_  (.A1(\heichips25_can_lehmann_fsm/net161 ),
    .A2(\heichips25_can_lehmann_fsm/_0535_ ),
    .Y(\heichips25_can_lehmann_fsm/_0036_ ),
    .B1(\heichips25_can_lehmann_fsm/_0536_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2208_  (.B1(\heichips25_can_lehmann_fsm/net1207 ),
    .Y(\heichips25_can_lehmann_fsm/_0537_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[9] ),
    .A2(\heichips25_can_lehmann_fsm/_1102_ ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_2209_  (.Y(\heichips25_can_lehmann_fsm/_0538_ ),
    .A(\heichips25_can_lehmann_fsm/_1103_ ),
    .B(\heichips25_can_lehmann_fsm/_0537_ ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_2210_  (.Y(\heichips25_can_lehmann_fsm/_0539_ ),
    .B1(\heichips25_can_lehmann_fsm/net165 ),
    .B2(\heichips25_can_lehmann_fsm/_0538_ ),
    .A2(\heichips25_can_lehmann_fsm/net176 ),
    .A1(\heichips25_can_lehmann_fsm/controller.const_data[10] ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2211_  (.B1(\heichips25_can_lehmann_fsm/net326 ),
    .Y(\heichips25_can_lehmann_fsm/_0540_ ),
    .A1(\heichips25_can_lehmann_fsm/net1207 ),
    .A2(\heichips25_can_lehmann_fsm/net161 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2212_  (.A1(\heichips25_can_lehmann_fsm/net161 ),
    .A2(\heichips25_can_lehmann_fsm/_0539_ ),
    .Y(\heichips25_can_lehmann_fsm/_0037_ ),
    .B1(\heichips25_can_lehmann_fsm/_0540_ ));
 sg13g2_xnor2_1 \heichips25_can_lehmann_fsm/_2213_  (.Y(\heichips25_can_lehmann_fsm/_0541_ ),
    .A(\heichips25_can_lehmann_fsm/net1186 ),
    .B(\heichips25_can_lehmann_fsm/_1103_ ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_2214_  (.Y(\heichips25_can_lehmann_fsm/_0542_ ),
    .B1(\heichips25_can_lehmann_fsm/net165 ),
    .B2(\heichips25_can_lehmann_fsm/_0541_ ),
    .A2(\heichips25_can_lehmann_fsm/net176 ),
    .A1(\heichips25_can_lehmann_fsm/net1006 ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2215_  (.B1(\heichips25_can_lehmann_fsm/net329 ),
    .Y(\heichips25_can_lehmann_fsm/_0543_ ),
    .A1(\heichips25_can_lehmann_fsm/net1186 ),
    .A2(\heichips25_can_lehmann_fsm/net162 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2216_  (.A1(\heichips25_can_lehmann_fsm/net162 ),
    .A2(\heichips25_can_lehmann_fsm/_0542_ ),
    .Y(\heichips25_can_lehmann_fsm/_0038_ ),
    .B1(\heichips25_can_lehmann_fsm/_0543_ ));
 sg13g2_xnor2_1 \heichips25_can_lehmann_fsm/_2217_  (.Y(\heichips25_can_lehmann_fsm/_0544_ ),
    .A(\heichips25_can_lehmann_fsm/net1231 ),
    .B(\heichips25_can_lehmann_fsm/_1104_ ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_2218_  (.Y(\heichips25_can_lehmann_fsm/_0545_ ),
    .B1(\heichips25_can_lehmann_fsm/net165 ),
    .B2(\heichips25_can_lehmann_fsm/_0544_ ),
    .A2(\heichips25_can_lehmann_fsm/net176 ),
    .A1(\heichips25_can_lehmann_fsm/net1034 ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2219_  (.B1(\heichips25_can_lehmann_fsm/net329 ),
    .Y(\heichips25_can_lehmann_fsm/_0546_ ),
    .A1(\heichips25_can_lehmann_fsm/net1231 ),
    .A2(\heichips25_can_lehmann_fsm/net162 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2220_  (.A1(\heichips25_can_lehmann_fsm/net162 ),
    .A2(\heichips25_can_lehmann_fsm/_0545_ ),
    .Y(\heichips25_can_lehmann_fsm/_0039_ ),
    .B1(\heichips25_can_lehmann_fsm/_0546_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2221_  (.B1(\heichips25_can_lehmann_fsm/net1217 ),
    .Y(\heichips25_can_lehmann_fsm/_0547_ ),
    .A1(\heichips25_can_lehmann_fsm/net1279 ),
    .A2(\heichips25_can_lehmann_fsm/_1104_ ));
 sg13g2_nand2b_1 \heichips25_can_lehmann_fsm/_2222_  (.Y(\heichips25_can_lehmann_fsm/_0548_ ),
    .B(\heichips25_can_lehmann_fsm/_0547_ ),
    .A_N(\heichips25_can_lehmann_fsm/_1105_ ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_2223_  (.Y(\heichips25_can_lehmann_fsm/_0549_ ),
    .B1(\heichips25_can_lehmann_fsm/net165 ),
    .B2(\heichips25_can_lehmann_fsm/_0548_ ),
    .A2(\heichips25_can_lehmann_fsm/net176 ),
    .A1(\heichips25_can_lehmann_fsm/net1050 ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2224_  (.B1(\heichips25_can_lehmann_fsm/net326 ),
    .Y(\heichips25_can_lehmann_fsm/_0550_ ),
    .A1(\heichips25_can_lehmann_fsm/net1217 ),
    .A2(\heichips25_can_lehmann_fsm/net161 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2225_  (.A1(\heichips25_can_lehmann_fsm/net161 ),
    .A2(\heichips25_can_lehmann_fsm/_0549_ ),
    .Y(\heichips25_can_lehmann_fsm/_0040_ ),
    .B1(\heichips25_can_lehmann_fsm/_0550_ ));
 sg13g2_xor2_1 \heichips25_can_lehmann_fsm/_2226_  (.B(\heichips25_can_lehmann_fsm/_1105_ ),
    .A(\heichips25_can_lehmann_fsm/net1221 ),
    .X(\heichips25_can_lehmann_fsm/_0551_ ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_2227_  (.Y(\heichips25_can_lehmann_fsm/_0552_ ),
    .B1(\heichips25_can_lehmann_fsm/net165 ),
    .B2(\heichips25_can_lehmann_fsm/_0551_ ),
    .A2(\heichips25_can_lehmann_fsm/net176 ),
    .A1(\heichips25_can_lehmann_fsm/net1115 ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2228_  (.B1(\heichips25_can_lehmann_fsm/net329 ),
    .Y(\heichips25_can_lehmann_fsm/_0553_ ),
    .A1(\heichips25_can_lehmann_fsm/net1221 ),
    .A2(\heichips25_can_lehmann_fsm/net162 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2229_  (.A1(\heichips25_can_lehmann_fsm/net162 ),
    .A2(\heichips25_can_lehmann_fsm/_0552_ ),
    .Y(\heichips25_can_lehmann_fsm/_0041_ ),
    .B1(\heichips25_can_lehmann_fsm/_0553_ ));
 sg13g2_xor2_1 \heichips25_can_lehmann_fsm/_2230_  (.B(\heichips25_can_lehmann_fsm/_1106_ ),
    .A(\heichips25_can_lehmann_fsm/net1205 ),
    .X(\heichips25_can_lehmann_fsm/_0554_ ));
 sg13g2_a22oi_1 \heichips25_can_lehmann_fsm/_2231_  (.Y(\heichips25_can_lehmann_fsm/_0555_ ),
    .B1(\heichips25_can_lehmann_fsm/_0496_ ),
    .B2(\heichips25_can_lehmann_fsm/_0554_ ),
    .A2(\heichips25_can_lehmann_fsm/net176 ),
    .A1(\heichips25_can_lehmann_fsm/net1002 ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2232_  (.B1(\heichips25_can_lehmann_fsm/net326 ),
    .Y(\heichips25_can_lehmann_fsm/_0556_ ),
    .A1(\heichips25_can_lehmann_fsm/net1205 ),
    .A2(\heichips25_can_lehmann_fsm/net161 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2233_  (.A1(\heichips25_can_lehmann_fsm/net161 ),
    .A2(\heichips25_can_lehmann_fsm/_0555_ ),
    .Y(\heichips25_can_lehmann_fsm/_0042_ ),
    .B1(\heichips25_can_lehmann_fsm/_0556_ ));
 sg13g2_nand2b_1 \heichips25_can_lehmann_fsm/_2234_  (.Y(\heichips25_can_lehmann_fsm/_0557_ ),
    .B(\heichips25_can_lehmann_fsm/_0492_ ),
    .A_N(\heichips25_can_lehmann_fsm/_0461_ ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_2235_  (.A(\heichips25_can_lehmann_fsm/net1212 ),
    .B(\heichips25_can_lehmann_fsm/net170 ),
    .Y(\heichips25_can_lehmann_fsm/_0558_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2236_  (.A1(\heichips25_can_lehmann_fsm/net857 ),
    .A2(\heichips25_can_lehmann_fsm/net170 ),
    .Y(\heichips25_can_lehmann_fsm/_0559_ ),
    .B1(\heichips25_can_lehmann_fsm/_0558_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2237_  (.B1(\heichips25_can_lehmann_fsm/net329 ),
    .Y(\heichips25_can_lehmann_fsm/_0560_ ),
    .A1(\heichips25_can_lehmann_fsm/net1212 ),
    .A2(\heichips25_can_lehmann_fsm/net205 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2238_  (.A1(\heichips25_can_lehmann_fsm/net205 ),
    .A2(\heichips25_can_lehmann_fsm/_0559_ ),
    .Y(\heichips25_can_lehmann_fsm/_0043_ ),
    .B1(\heichips25_can_lehmann_fsm/_0560_ ));
 sg13g2_xor2_1 \heichips25_can_lehmann_fsm/_2239_  (.B(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[0] ),
    .A(\heichips25_can_lehmann_fsm/net1174 ),
    .X(\heichips25_can_lehmann_fsm/_0561_ ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_2240_  (.A(\heichips25_can_lehmann_fsm/net170 ),
    .B(\heichips25_can_lehmann_fsm/_0561_ ),
    .Y(\heichips25_can_lehmann_fsm/_0562_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2241_  (.A1(\heichips25_can_lehmann_fsm/net840 ),
    .A2(\heichips25_can_lehmann_fsm/net170 ),
    .Y(\heichips25_can_lehmann_fsm/_0563_ ),
    .B1(\heichips25_can_lehmann_fsm/_0562_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2242_  (.B1(\heichips25_can_lehmann_fsm/net329 ),
    .Y(\heichips25_can_lehmann_fsm/_0564_ ),
    .A1(\heichips25_can_lehmann_fsm/net1174 ),
    .A2(\heichips25_can_lehmann_fsm/net205 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2243_  (.A1(\heichips25_can_lehmann_fsm/net205 ),
    .A2(\heichips25_can_lehmann_fsm/_0563_ ),
    .Y(\heichips25_can_lehmann_fsm/_0044_ ),
    .B1(\heichips25_can_lehmann_fsm/_0564_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2244_  (.B1(\heichips25_can_lehmann_fsm/net1195 ),
    .Y(\heichips25_can_lehmann_fsm/_0565_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[1] ),
    .A2(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[0] ));
 sg13g2_nor2b_1 \heichips25_can_lehmann_fsm/_2245_  (.A(\heichips25_can_lehmann_fsm/_1043_ ),
    .B_N(\heichips25_can_lehmann_fsm/_0565_ ),
    .Y(\heichips25_can_lehmann_fsm/_0566_ ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_2246_  (.A(\heichips25_can_lehmann_fsm/net170 ),
    .B(\heichips25_can_lehmann_fsm/_0566_ ),
    .Y(\heichips25_can_lehmann_fsm/_0567_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2247_  (.A1(\heichips25_can_lehmann_fsm/net911 ),
    .A2(\heichips25_can_lehmann_fsm/net170 ),
    .Y(\heichips25_can_lehmann_fsm/_0568_ ),
    .B1(\heichips25_can_lehmann_fsm/_0567_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2248_  (.B1(\heichips25_can_lehmann_fsm/net329 ),
    .Y(\heichips25_can_lehmann_fsm/_0569_ ),
    .A1(\heichips25_can_lehmann_fsm/net1195 ),
    .A2(\heichips25_can_lehmann_fsm/net210 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2249_  (.A1(\heichips25_can_lehmann_fsm/net210 ),
    .A2(\heichips25_can_lehmann_fsm/_0568_ ),
    .Y(\heichips25_can_lehmann_fsm/_0045_ ),
    .B1(\heichips25_can_lehmann_fsm/_0569_ ));
 sg13g2_nand2b_1 \heichips25_can_lehmann_fsm/_2250_  (.Y(\heichips25_can_lehmann_fsm/_0570_ ),
    .B(\heichips25_can_lehmann_fsm/net1173 ),
    .A_N(\heichips25_can_lehmann_fsm/_1043_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2251_  (.A1(\heichips25_can_lehmann_fsm/_1044_ ),
    .A2(\heichips25_can_lehmann_fsm/_0570_ ),
    .Y(\heichips25_can_lehmann_fsm/_0571_ ),
    .B1(\heichips25_can_lehmann_fsm/net170 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2252_  (.A1(\heichips25_can_lehmann_fsm/net898 ),
    .A2(\heichips25_can_lehmann_fsm/net170 ),
    .Y(\heichips25_can_lehmann_fsm/_0572_ ),
    .B1(\heichips25_can_lehmann_fsm/_0571_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2253_  (.B1(\heichips25_can_lehmann_fsm/net327 ),
    .Y(\heichips25_can_lehmann_fsm/_0573_ ),
    .A1(\heichips25_can_lehmann_fsm/net1173 ),
    .A2(\heichips25_can_lehmann_fsm/net206 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2254_  (.A1(\heichips25_can_lehmann_fsm/net206 ),
    .A2(\heichips25_can_lehmann_fsm/_0572_ ),
    .Y(\heichips25_can_lehmann_fsm/_0046_ ),
    .B1(\heichips25_can_lehmann_fsm/_0573_ ));
 sg13g2_xor2_1 \heichips25_can_lehmann_fsm/_2255_  (.B(\heichips25_can_lehmann_fsm/_1044_ ),
    .A(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[4] ),
    .X(\heichips25_can_lehmann_fsm/_0574_ ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_2256_  (.A(\heichips25_can_lehmann_fsm/net173 ),
    .B(\heichips25_can_lehmann_fsm/_0574_ ),
    .Y(\heichips25_can_lehmann_fsm/_0575_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2257_  (.A1(\heichips25_can_lehmann_fsm/net1183 ),
    .A2(\heichips25_can_lehmann_fsm/net173 ),
    .Y(\heichips25_can_lehmann_fsm/_0576_ ),
    .B1(\heichips25_can_lehmann_fsm/_0575_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2258_  (.B1(\heichips25_can_lehmann_fsm/net327 ),
    .Y(\heichips25_can_lehmann_fsm/_0577_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[4] ),
    .A2(\heichips25_can_lehmann_fsm/net206 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2259_  (.A1(\heichips25_can_lehmann_fsm/net206 ),
    .A2(\heichips25_can_lehmann_fsm/net1184 ),
    .Y(\heichips25_can_lehmann_fsm/_0047_ ),
    .B1(\heichips25_can_lehmann_fsm/_0577_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2260_  (.B1(\heichips25_can_lehmann_fsm/net1181 ),
    .Y(\heichips25_can_lehmann_fsm/_0578_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[4] ),
    .A2(\heichips25_can_lehmann_fsm/_1044_ ));
 sg13g2_nor2b_1 \heichips25_can_lehmann_fsm/_2261_  (.A(\heichips25_can_lehmann_fsm/_1045_ ),
    .B_N(\heichips25_can_lehmann_fsm/_0578_ ),
    .Y(\heichips25_can_lehmann_fsm/_0579_ ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_2262_  (.A(\heichips25_can_lehmann_fsm/net173 ),
    .B(\heichips25_can_lehmann_fsm/_0579_ ),
    .Y(\heichips25_can_lehmann_fsm/_0580_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2263_  (.A1(\heichips25_can_lehmann_fsm/net939 ),
    .A2(\heichips25_can_lehmann_fsm/net173 ),
    .Y(\heichips25_can_lehmann_fsm/_0581_ ),
    .B1(\heichips25_can_lehmann_fsm/_0580_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2264_  (.B1(\heichips25_can_lehmann_fsm/net327 ),
    .Y(\heichips25_can_lehmann_fsm/_0582_ ),
    .A1(\heichips25_can_lehmann_fsm/net1181 ),
    .A2(\heichips25_can_lehmann_fsm/net208 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2265_  (.A1(\heichips25_can_lehmann_fsm/net208 ),
    .A2(\heichips25_can_lehmann_fsm/_0581_ ),
    .Y(\heichips25_can_lehmann_fsm/_0048_ ),
    .B1(\heichips25_can_lehmann_fsm/_0582_ ));
 sg13g2_xnor2_1 \heichips25_can_lehmann_fsm/_2266_  (.Y(\heichips25_can_lehmann_fsm/_0583_ ),
    .A(\heichips25_can_lehmann_fsm/net1194 ),
    .B(\heichips25_can_lehmann_fsm/_1045_ ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_2267_  (.A(\heichips25_can_lehmann_fsm/net171 ),
    .B(\heichips25_can_lehmann_fsm/_0583_ ),
    .Y(\heichips25_can_lehmann_fsm/_0584_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2268_  (.A1(\heichips25_can_lehmann_fsm/net941 ),
    .A2(\heichips25_can_lehmann_fsm/net171 ),
    .Y(\heichips25_can_lehmann_fsm/_0585_ ),
    .B1(\heichips25_can_lehmann_fsm/_0584_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2269_  (.B1(\heichips25_can_lehmann_fsm/net327 ),
    .Y(\heichips25_can_lehmann_fsm/_0586_ ),
    .A1(\heichips25_can_lehmann_fsm/net1194 ),
    .A2(\heichips25_can_lehmann_fsm/net207 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2270_  (.A1(\heichips25_can_lehmann_fsm/net207 ),
    .A2(\heichips25_can_lehmann_fsm/_0585_ ),
    .Y(\heichips25_can_lehmann_fsm/_0049_ ),
    .B1(\heichips25_can_lehmann_fsm/_0586_ ));
 sg13g2_nand2b_1 \heichips25_can_lehmann_fsm/_2271_  (.Y(\heichips25_can_lehmann_fsm/_0587_ ),
    .B(\heichips25_can_lehmann_fsm/net1182 ),
    .A_N(\heichips25_can_lehmann_fsm/_1046_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2272_  (.A1(\heichips25_can_lehmann_fsm/_1047_ ),
    .A2(\heichips25_can_lehmann_fsm/_0587_ ),
    .Y(\heichips25_can_lehmann_fsm/_0588_ ),
    .B1(\heichips25_can_lehmann_fsm/net172 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2273_  (.A1(\heichips25_can_lehmann_fsm/net965 ),
    .A2(\heichips25_can_lehmann_fsm/net172 ),
    .Y(\heichips25_can_lehmann_fsm/_0589_ ),
    .B1(\heichips25_can_lehmann_fsm/_0588_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2274_  (.B1(\heichips25_can_lehmann_fsm/net327 ),
    .Y(\heichips25_can_lehmann_fsm/_0590_ ),
    .A1(\heichips25_can_lehmann_fsm/net1182 ),
    .A2(\heichips25_can_lehmann_fsm/net207 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2275_  (.A1(\heichips25_can_lehmann_fsm/net207 ),
    .A2(\heichips25_can_lehmann_fsm/_0589_ ),
    .Y(\heichips25_can_lehmann_fsm/_0050_ ),
    .B1(\heichips25_can_lehmann_fsm/_0590_ ));
 sg13g2_xor2_1 \heichips25_can_lehmann_fsm/_2276_  (.B(\heichips25_can_lehmann_fsm/_1047_ ),
    .A(\heichips25_can_lehmann_fsm/net1191 ),
    .X(\heichips25_can_lehmann_fsm/_0591_ ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_2277_  (.A(\heichips25_can_lehmann_fsm/net172 ),
    .B(\heichips25_can_lehmann_fsm/_0591_ ),
    .Y(\heichips25_can_lehmann_fsm/_0592_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2278_  (.A1(\heichips25_can_lehmann_fsm/net968 ),
    .A2(\heichips25_can_lehmann_fsm/net172 ),
    .Y(\heichips25_can_lehmann_fsm/_0593_ ),
    .B1(\heichips25_can_lehmann_fsm/_0592_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2279_  (.B1(\heichips25_can_lehmann_fsm/net328 ),
    .Y(\heichips25_can_lehmann_fsm/_0594_ ),
    .A1(\heichips25_can_lehmann_fsm/net1191 ),
    .A2(\heichips25_can_lehmann_fsm/net208 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2280_  (.A1(\heichips25_can_lehmann_fsm/net208 ),
    .A2(\heichips25_can_lehmann_fsm/_0593_ ),
    .Y(\heichips25_can_lehmann_fsm/_0051_ ),
    .B1(\heichips25_can_lehmann_fsm/_0594_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2281_  (.B1(\heichips25_can_lehmann_fsm/net1170 ),
    .Y(\heichips25_can_lehmann_fsm/_0595_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[8] ),
    .A2(\heichips25_can_lehmann_fsm/_1047_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2282_  (.A1(\heichips25_can_lehmann_fsm/_1049_ ),
    .A2(\heichips25_can_lehmann_fsm/_0595_ ),
    .Y(\heichips25_can_lehmann_fsm/_0596_ ),
    .B1(\heichips25_can_lehmann_fsm/net171 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2283_  (.A1(\heichips25_can_lehmann_fsm/net942 ),
    .A2(\heichips25_can_lehmann_fsm/net171 ),
    .Y(\heichips25_can_lehmann_fsm/_0597_ ),
    .B1(\heichips25_can_lehmann_fsm/_0596_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2284_  (.B1(\heichips25_can_lehmann_fsm/net328 ),
    .Y(\heichips25_can_lehmann_fsm/_0598_ ),
    .A1(\heichips25_can_lehmann_fsm/net1170 ),
    .A2(\heichips25_can_lehmann_fsm/net207 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2285_  (.A1(\heichips25_can_lehmann_fsm/net207 ),
    .A2(\heichips25_can_lehmann_fsm/_0597_ ),
    .Y(\heichips25_can_lehmann_fsm/_0052_ ),
    .B1(\heichips25_can_lehmann_fsm/_0598_ ));
 sg13g2_xor2_1 \heichips25_can_lehmann_fsm/_2286_  (.B(\heichips25_can_lehmann_fsm/_1049_ ),
    .A(\heichips25_can_lehmann_fsm/net1209 ),
    .X(\heichips25_can_lehmann_fsm/_0599_ ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_2287_  (.A(\heichips25_can_lehmann_fsm/net171 ),
    .B(\heichips25_can_lehmann_fsm/_0599_ ),
    .Y(\heichips25_can_lehmann_fsm/_0600_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2288_  (.A1(\heichips25_can_lehmann_fsm/net980 ),
    .A2(\heichips25_can_lehmann_fsm/net171 ),
    .Y(\heichips25_can_lehmann_fsm/_0601_ ),
    .B1(\heichips25_can_lehmann_fsm/_0600_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2289_  (.B1(\heichips25_can_lehmann_fsm/net328 ),
    .Y(\heichips25_can_lehmann_fsm/_0602_ ),
    .A1(\heichips25_can_lehmann_fsm/net1209 ),
    .A2(\heichips25_can_lehmann_fsm/net207 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2290_  (.A1(\heichips25_can_lehmann_fsm/net207 ),
    .A2(\heichips25_can_lehmann_fsm/_0601_ ),
    .Y(\heichips25_can_lehmann_fsm/_0053_ ),
    .B1(\heichips25_can_lehmann_fsm/_0602_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2291_  (.B1(\heichips25_can_lehmann_fsm/net1165 ),
    .Y(\heichips25_can_lehmann_fsm/_0603_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[10] ),
    .A2(\heichips25_can_lehmann_fsm/_1049_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2292_  (.A1(\heichips25_can_lehmann_fsm/_1051_ ),
    .A2(\heichips25_can_lehmann_fsm/_0603_ ),
    .Y(\heichips25_can_lehmann_fsm/_0604_ ),
    .B1(\heichips25_can_lehmann_fsm/net171 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2293_  (.A1(\heichips25_can_lehmann_fsm/net948 ),
    .A2(\heichips25_can_lehmann_fsm/net171 ),
    .Y(\heichips25_can_lehmann_fsm/_0605_ ),
    .B1(\heichips25_can_lehmann_fsm/_0604_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2294_  (.B1(\heichips25_can_lehmann_fsm/net328 ),
    .Y(\heichips25_can_lehmann_fsm/_0606_ ),
    .A1(\heichips25_can_lehmann_fsm/net1165 ),
    .A2(\heichips25_can_lehmann_fsm/net208 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2295_  (.A1(\heichips25_can_lehmann_fsm/net208 ),
    .A2(\heichips25_can_lehmann_fsm/_0605_ ),
    .Y(\heichips25_can_lehmann_fsm/_0054_ ),
    .B1(\heichips25_can_lehmann_fsm/_0606_ ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_2296_  (.Y(\heichips25_can_lehmann_fsm/_0607_ ),
    .A(\heichips25_can_lehmann_fsm/net206 ),
    .B(\heichips25_can_lehmann_fsm/net174 ));
 sg13g2_nor2b_1 \heichips25_can_lehmann_fsm/_2297_  (.A(\heichips25_can_lehmann_fsm/_1051_ ),
    .B_N(\heichips25_can_lehmann_fsm/net209 ),
    .Y(\heichips25_can_lehmann_fsm/_0608_ ));
 sg13g2_xnor2_1 \heichips25_can_lehmann_fsm/_2298_  (.Y(\heichips25_can_lehmann_fsm/_0609_ ),
    .A(\heichips25_can_lehmann_fsm/net1200 ),
    .B(\heichips25_can_lehmann_fsm/_0608_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2299_  (.B1(\heichips25_can_lehmann_fsm/net327 ),
    .Y(\heichips25_can_lehmann_fsm/_0610_ ),
    .A1(\heichips25_can_lehmann_fsm/net983 ),
    .A2(\heichips25_can_lehmann_fsm/_0607_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2300_  (.A1(\heichips25_can_lehmann_fsm/_0607_ ),
    .A2(\heichips25_can_lehmann_fsm/net1201 ),
    .Y(\heichips25_can_lehmann_fsm/_0055_ ),
    .B1(\heichips25_can_lehmann_fsm/_0610_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2301_  (.B1(\heichips25_can_lehmann_fsm/net1158 ),
    .Y(\heichips25_can_lehmann_fsm/_0611_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[12] ),
    .A2(\heichips25_can_lehmann_fsm/_1051_ ));
 sg13g2_nor2b_1 \heichips25_can_lehmann_fsm/_2302_  (.A(\heichips25_can_lehmann_fsm/_1052_ ),
    .B_N(\heichips25_can_lehmann_fsm/_0611_ ),
    .Y(\heichips25_can_lehmann_fsm/_0612_ ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_2303_  (.A(\heichips25_can_lehmann_fsm/net173 ),
    .B(\heichips25_can_lehmann_fsm/_0612_ ),
    .Y(\heichips25_can_lehmann_fsm/_0613_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2304_  (.A1(\heichips25_can_lehmann_fsm/net1085 ),
    .A2(\heichips25_can_lehmann_fsm/net173 ),
    .Y(\heichips25_can_lehmann_fsm/_0614_ ),
    .B1(\heichips25_can_lehmann_fsm/_0613_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2305_  (.B1(\heichips25_can_lehmann_fsm/net327 ),
    .Y(\heichips25_can_lehmann_fsm/_0615_ ),
    .A1(\heichips25_can_lehmann_fsm/net1158 ),
    .A2(\heichips25_can_lehmann_fsm/net209 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2306_  (.A1(\heichips25_can_lehmann_fsm/net209 ),
    .A2(\heichips25_can_lehmann_fsm/_0614_ ),
    .Y(\heichips25_can_lehmann_fsm/_0056_ ),
    .B1(\heichips25_can_lehmann_fsm/_0615_ ));
 sg13g2_xnor2_1 \heichips25_can_lehmann_fsm/_2307_  (.Y(\heichips25_can_lehmann_fsm/_0616_ ),
    .A(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[14] ),
    .B(\heichips25_can_lehmann_fsm/_1052_ ));
 sg13g2_nor2_1 \heichips25_can_lehmann_fsm/_2308_  (.A(\heichips25_can_lehmann_fsm/net174 ),
    .B(\heichips25_can_lehmann_fsm/_0616_ ),
    .Y(\heichips25_can_lehmann_fsm/_0617_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2309_  (.A1(\heichips25_can_lehmann_fsm/net1188 ),
    .A2(\heichips25_can_lehmann_fsm/net174 ),
    .Y(\heichips25_can_lehmann_fsm/_0618_ ),
    .B1(\heichips25_can_lehmann_fsm/_0617_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2310_  (.B1(\heichips25_can_lehmann_fsm/net327 ),
    .Y(\heichips25_can_lehmann_fsm/_0619_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[14] ),
    .A2(\heichips25_can_lehmann_fsm/net206 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2311_  (.A1(\heichips25_can_lehmann_fsm/net206 ),
    .A2(\heichips25_can_lehmann_fsm/net1189 ),
    .Y(\heichips25_can_lehmann_fsm/_0057_ ),
    .B1(\heichips25_can_lehmann_fsm/_0619_ ));
 sg13g2_nand3b_1 \heichips25_can_lehmann_fsm/_2312_  (.B(\heichips25_can_lehmann_fsm/_1052_ ),
    .C(\heichips25_can_lehmann_fsm/net206 ),
    .Y(\heichips25_can_lehmann_fsm/_0620_ ),
    .A_N(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[14] ));
 sg13g2_xor2_1 \heichips25_can_lehmann_fsm/_2313_  (.B(\heichips25_can_lehmann_fsm/_0620_ ),
    .A(\heichips25_can_lehmann_fsm/net1168 ),
    .X(\heichips25_can_lehmann_fsm/_0621_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2314_  (.B1(\heichips25_can_lehmann_fsm/net329 ),
    .Y(\heichips25_can_lehmann_fsm/_0622_ ),
    .A1(\heichips25_can_lehmann_fsm/net883 ),
    .A2(\heichips25_can_lehmann_fsm/_0607_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2315_  (.A1(\heichips25_can_lehmann_fsm/_0607_ ),
    .A2(\heichips25_can_lehmann_fsm/net1169 ),
    .Y(\heichips25_can_lehmann_fsm/_0058_ ),
    .B1(\heichips25_can_lehmann_fsm/_0622_ ));
 sg13g2_and2_1 \heichips25_can_lehmann_fsm/_2316_  (.A(net8),
    .B(net9),
    .X(\heichips25_can_lehmann_fsm/_0623_ ));
 sg13g2_nand2_1 \heichips25_can_lehmann_fsm/_2317_  (.Y(\heichips25_can_lehmann_fsm/_0624_ ),
    .A(net8),
    .B(net9));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2318_  (.B1(\heichips25_can_lehmann_fsm/net473 ),
    .Y(\heichips25_can_lehmann_fsm/_0625_ ),
    .A1(\heichips25_can_lehmann_fsm/net1204 ),
    .A2(\heichips25_can_lehmann_fsm/net401 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2319_  (.A1(\heichips25_can_lehmann_fsm/_0972_ ),
    .A2(\heichips25_can_lehmann_fsm/net401 ),
    .Y(\heichips25_can_lehmann_fsm/_0059_ ),
    .B1(\heichips25_can_lehmann_fsm/_0625_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2320_  (.B1(\heichips25_can_lehmann_fsm/net474 ),
    .Y(\heichips25_can_lehmann_fsm/_0626_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.const_data[0] ),
    .A2(\heichips25_can_lehmann_fsm/net363 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2321_  (.A1(\heichips25_can_lehmann_fsm/_0971_ ),
    .A2(\heichips25_can_lehmann_fsm/net363 ),
    .Y(\heichips25_can_lehmann_fsm/_0060_ ),
    .B1(\heichips25_can_lehmann_fsm/_0626_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2322_  (.B1(\heichips25_can_lehmann_fsm/net471 ),
    .Y(\heichips25_can_lehmann_fsm/_0627_ ),
    .A1(\heichips25_can_lehmann_fsm/net1136 ),
    .A2(\heichips25_can_lehmann_fsm/net403 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2323_  (.A1(\heichips25_can_lehmann_fsm/_0971_ ),
    .A2(\heichips25_can_lehmann_fsm/net403 ),
    .Y(\heichips25_can_lehmann_fsm/_0061_ ),
    .B1(\heichips25_can_lehmann_fsm/_0627_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2324_  (.B1(\heichips25_can_lehmann_fsm/net471 ),
    .Y(\heichips25_can_lehmann_fsm/_0628_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.const_data[2] ),
    .A2(\heichips25_can_lehmann_fsm/net363 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2325_  (.A1(\heichips25_can_lehmann_fsm/_0970_ ),
    .A2(\heichips25_can_lehmann_fsm/net363 ),
    .Y(\heichips25_can_lehmann_fsm/_0062_ ),
    .B1(\heichips25_can_lehmann_fsm/_0628_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2326_  (.B1(\heichips25_can_lehmann_fsm/net471 ),
    .Y(\heichips25_can_lehmann_fsm/_0629_ ),
    .A1(\heichips25_can_lehmann_fsm/net933 ),
    .A2(\heichips25_can_lehmann_fsm/net403 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2327_  (.A1(\heichips25_can_lehmann_fsm/_0970_ ),
    .A2(\heichips25_can_lehmann_fsm/net403 ),
    .Y(\heichips25_can_lehmann_fsm/_0063_ ),
    .B1(\heichips25_can_lehmann_fsm/_0629_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2328_  (.B1(\heichips25_can_lehmann_fsm/net471 ),
    .Y(\heichips25_can_lehmann_fsm/_0630_ ),
    .A1(\heichips25_can_lehmann_fsm/net933 ),
    .A2(\heichips25_can_lehmann_fsm/net363 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2329_  (.A1(\heichips25_can_lehmann_fsm/_0969_ ),
    .A2(\heichips25_can_lehmann_fsm/net363 ),
    .Y(\heichips25_can_lehmann_fsm/_0064_ ),
    .B1(\heichips25_can_lehmann_fsm/_0630_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2330_  (.B1(\heichips25_can_lehmann_fsm/net471 ),
    .Y(\heichips25_can_lehmann_fsm/_0631_ ),
    .A1(\heichips25_can_lehmann_fsm/net1113 ),
    .A2(\heichips25_can_lehmann_fsm/net403 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2331_  (.A1(\heichips25_can_lehmann_fsm/_0969_ ),
    .A2(\heichips25_can_lehmann_fsm/net403 ),
    .Y(\heichips25_can_lehmann_fsm/_0065_ ),
    .B1(\heichips25_can_lehmann_fsm/_0631_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2332_  (.B1(\heichips25_can_lehmann_fsm/net475 ),
    .Y(\heichips25_can_lehmann_fsm/_0632_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.const_data[6] ),
    .A2(\heichips25_can_lehmann_fsm/net363 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2333_  (.A1(\heichips25_can_lehmann_fsm/_0968_ ),
    .A2(\heichips25_can_lehmann_fsm/net363 ),
    .Y(\heichips25_can_lehmann_fsm/_0066_ ),
    .B1(\heichips25_can_lehmann_fsm/_0632_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2334_  (.B1(\heichips25_can_lehmann_fsm/net474 ),
    .Y(\heichips25_can_lehmann_fsm/_0633_ ),
    .A1(\heichips25_can_lehmann_fsm/net974 ),
    .A2(\heichips25_can_lehmann_fsm/net403 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2335_  (.A1(\heichips25_can_lehmann_fsm/_0968_ ),
    .A2(\heichips25_can_lehmann_fsm/net408 ),
    .Y(\heichips25_can_lehmann_fsm/_0067_ ),
    .B1(\heichips25_can_lehmann_fsm/_0633_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2336_  (.B1(\heichips25_can_lehmann_fsm/net474 ),
    .Y(\heichips25_can_lehmann_fsm/_0634_ ),
    .A1(\heichips25_can_lehmann_fsm/net974 ),
    .A2(\heichips25_can_lehmann_fsm/net364 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2337_  (.A1(\heichips25_can_lehmann_fsm/_0967_ ),
    .A2(\heichips25_can_lehmann_fsm/net367 ),
    .Y(\heichips25_can_lehmann_fsm/_0068_ ),
    .B1(\heichips25_can_lehmann_fsm/_0634_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2338_  (.B1(\heichips25_can_lehmann_fsm/net474 ),
    .Y(\heichips25_can_lehmann_fsm/_0635_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.const_data[10] ),
    .A2(\heichips25_can_lehmann_fsm/net406 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2339_  (.A1(\heichips25_can_lehmann_fsm/_0967_ ),
    .A2(\heichips25_can_lehmann_fsm/net406 ),
    .Y(\heichips25_can_lehmann_fsm/_0069_ ),
    .B1(\heichips25_can_lehmann_fsm/_0635_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2340_  (.B1(\heichips25_can_lehmann_fsm/net474 ),
    .Y(\heichips25_can_lehmann_fsm/_0636_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.const_data[10] ),
    .A2(\heichips25_can_lehmann_fsm/net367 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2341_  (.A1(\heichips25_can_lehmann_fsm/_0966_ ),
    .A2(\heichips25_can_lehmann_fsm/net367 ),
    .Y(\heichips25_can_lehmann_fsm/_0070_ ),
    .B1(\heichips25_can_lehmann_fsm/_0636_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2342_  (.B1(\heichips25_can_lehmann_fsm/net494 ),
    .Y(\heichips25_can_lehmann_fsm/_0637_ ),
    .A1(\heichips25_can_lehmann_fsm/net1034 ),
    .A2(\heichips25_can_lehmann_fsm/net406 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2343_  (.A1(\heichips25_can_lehmann_fsm/_0966_ ),
    .A2(\heichips25_can_lehmann_fsm/net406 ),
    .Y(\heichips25_can_lehmann_fsm/_0071_ ),
    .B1(\heichips25_can_lehmann_fsm/_0637_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2344_  (.B1(\heichips25_can_lehmann_fsm/net494 ),
    .Y(\heichips25_can_lehmann_fsm/_0638_ ),
    .A1(\heichips25_can_lehmann_fsm/net1034 ),
    .A2(\heichips25_can_lehmann_fsm/net367 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2345_  (.A1(\heichips25_can_lehmann_fsm/_0965_ ),
    .A2(\heichips25_can_lehmann_fsm/net367 ),
    .Y(\heichips25_can_lehmann_fsm/_0072_ ),
    .B1(\heichips25_can_lehmann_fsm/_0638_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2346_  (.B1(\heichips25_can_lehmann_fsm/net494 ),
    .Y(\heichips25_can_lehmann_fsm/_0639_ ),
    .A1(\heichips25_can_lehmann_fsm/net1115 ),
    .A2(\heichips25_can_lehmann_fsm/net406 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2347_  (.A1(\heichips25_can_lehmann_fsm/_0965_ ),
    .A2(\heichips25_can_lehmann_fsm/net406 ),
    .Y(\heichips25_can_lehmann_fsm/_0073_ ),
    .B1(\heichips25_can_lehmann_fsm/_0639_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2348_  (.B1(\heichips25_can_lehmann_fsm/net494 ),
    .Y(\heichips25_can_lehmann_fsm/_0640_ ),
    .A1(\heichips25_can_lehmann_fsm/net1115 ),
    .A2(\heichips25_can_lehmann_fsm/net382 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2349_  (.A1(\heichips25_can_lehmann_fsm/_0964_ ),
    .A2(\heichips25_can_lehmann_fsm/net382 ),
    .Y(\heichips25_can_lehmann_fsm/_0074_ ),
    .B1(\heichips25_can_lehmann_fsm/_0640_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2350_  (.B1(\heichips25_can_lehmann_fsm/net494 ),
    .Y(\heichips25_can_lehmann_fsm/_0641_ ),
    .A1(\heichips25_can_lehmann_fsm/net857 ),
    .A2(\heichips25_can_lehmann_fsm/net423 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2351_  (.A1(\heichips25_can_lehmann_fsm/_0964_ ),
    .A2(\heichips25_can_lehmann_fsm/net423 ),
    .Y(\heichips25_can_lehmann_fsm/_0075_ ),
    .B1(\heichips25_can_lehmann_fsm/_0641_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2352_  (.B1(\heichips25_can_lehmann_fsm/net494 ),
    .Y(\heichips25_can_lehmann_fsm/_0642_ ),
    .A1(\heichips25_can_lehmann_fsm/net857 ),
    .A2(\heichips25_can_lehmann_fsm/net383 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2353_  (.A1(\heichips25_can_lehmann_fsm/_0963_ ),
    .A2(\heichips25_can_lehmann_fsm/net383 ),
    .Y(\heichips25_can_lehmann_fsm/_0076_ ),
    .B1(\heichips25_can_lehmann_fsm/_0642_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2354_  (.B1(\heichips25_can_lehmann_fsm/net495 ),
    .Y(\heichips25_can_lehmann_fsm/_0643_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.const_data[18] ),
    .A2(\heichips25_can_lehmann_fsm/net423 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2355_  (.A1(\heichips25_can_lehmann_fsm/_0963_ ),
    .A2(\heichips25_can_lehmann_fsm/net423 ),
    .Y(\heichips25_can_lehmann_fsm/_0077_ ),
    .B1(\heichips25_can_lehmann_fsm/_0643_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2356_  (.B1(\heichips25_can_lehmann_fsm/net495 ),
    .Y(\heichips25_can_lehmann_fsm/_0644_ ),
    .A1(\heichips25_can_lehmann_fsm/net911 ),
    .A2(\heichips25_can_lehmann_fsm/net383 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2357_  (.A1(\heichips25_can_lehmann_fsm/_0962_ ),
    .A2(\heichips25_can_lehmann_fsm/net383 ),
    .Y(\heichips25_can_lehmann_fsm/_0078_ ),
    .B1(\heichips25_can_lehmann_fsm/_0644_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2358_  (.B1(\heichips25_can_lehmann_fsm/net500 ),
    .Y(\heichips25_can_lehmann_fsm/_0645_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.const_data[20] ),
    .A2(\heichips25_can_lehmann_fsm/net424 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2359_  (.A1(\heichips25_can_lehmann_fsm/_0962_ ),
    .A2(\heichips25_can_lehmann_fsm/net424 ),
    .Y(\heichips25_can_lehmann_fsm/_0079_ ),
    .B1(\heichips25_can_lehmann_fsm/_0645_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2360_  (.B1(\heichips25_can_lehmann_fsm/net500 ),
    .Y(\heichips25_can_lehmann_fsm/_0646_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.const_data[20] ),
    .A2(\heichips25_can_lehmann_fsm/net387 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2361_  (.A1(\heichips25_can_lehmann_fsm/_0961_ ),
    .A2(\heichips25_can_lehmann_fsm/net387 ),
    .Y(\heichips25_can_lehmann_fsm/_0080_ ),
    .B1(\heichips25_can_lehmann_fsm/_0646_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2362_  (.B1(\heichips25_can_lehmann_fsm/net500 ),
    .Y(\heichips25_can_lehmann_fsm/_0647_ ),
    .A1(\heichips25_can_lehmann_fsm/net941 ),
    .A2(\heichips25_can_lehmann_fsm/net430 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2363_  (.A1(\heichips25_can_lehmann_fsm/_0961_ ),
    .A2(\heichips25_can_lehmann_fsm/net430 ),
    .Y(\heichips25_can_lehmann_fsm/_0081_ ),
    .B1(\heichips25_can_lehmann_fsm/_0647_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2364_  (.B1(\heichips25_can_lehmann_fsm/net500 ),
    .Y(\heichips25_can_lehmann_fsm/_0648_ ),
    .A1(\heichips25_can_lehmann_fsm/net941 ),
    .A2(\heichips25_can_lehmann_fsm/net387 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2365_  (.A1(\heichips25_can_lehmann_fsm/_0960_ ),
    .A2(\heichips25_can_lehmann_fsm/net387 ),
    .Y(\heichips25_can_lehmann_fsm/_0082_ ),
    .B1(\heichips25_can_lehmann_fsm/_0648_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2366_  (.B1(\heichips25_can_lehmann_fsm/net501 ),
    .Y(\heichips25_can_lehmann_fsm/_0649_ ),
    .A1(\heichips25_can_lehmann_fsm/net968 ),
    .A2(\heichips25_can_lehmann_fsm/net430 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2367_  (.A1(\heichips25_can_lehmann_fsm/_0960_ ),
    .A2(\heichips25_can_lehmann_fsm/net431 ),
    .Y(\heichips25_can_lehmann_fsm/_0083_ ),
    .B1(\heichips25_can_lehmann_fsm/_0649_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2368_  (.B1(\heichips25_can_lehmann_fsm/net501 ),
    .Y(\heichips25_can_lehmann_fsm/_0650_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.const_data[24] ),
    .A2(\heichips25_can_lehmann_fsm/net387 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2369_  (.A1(\heichips25_can_lehmann_fsm/_0959_ ),
    .A2(\heichips25_can_lehmann_fsm/net388 ),
    .Y(\heichips25_can_lehmann_fsm/_0084_ ),
    .B1(\heichips25_can_lehmann_fsm/_0650_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2370_  (.B1(\heichips25_can_lehmann_fsm/net501 ),
    .Y(\heichips25_can_lehmann_fsm/_0651_ ),
    .A1(\heichips25_can_lehmann_fsm/net980 ),
    .A2(\heichips25_can_lehmann_fsm/net431 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2371_  (.A1(\heichips25_can_lehmann_fsm/_0959_ ),
    .A2(\heichips25_can_lehmann_fsm/net431 ),
    .Y(\heichips25_can_lehmann_fsm/_0085_ ),
    .B1(\heichips25_can_lehmann_fsm/_0651_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2372_  (.B1(\heichips25_can_lehmann_fsm/net501 ),
    .Y(\heichips25_can_lehmann_fsm/_0652_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.const_data[26] ),
    .A2(\heichips25_can_lehmann_fsm/net388 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2373_  (.A1(\heichips25_can_lehmann_fsm/_0958_ ),
    .A2(\heichips25_can_lehmann_fsm/net388 ),
    .Y(\heichips25_can_lehmann_fsm/_0086_ ),
    .B1(\heichips25_can_lehmann_fsm/_0652_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2374_  (.B1(\heichips25_can_lehmann_fsm/net500 ),
    .Y(\heichips25_can_lehmann_fsm/_0653_ ),
    .A1(\heichips25_can_lehmann_fsm/net983 ),
    .A2(\heichips25_can_lehmann_fsm/net430 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2375_  (.A1(\heichips25_can_lehmann_fsm/_0958_ ),
    .A2(\heichips25_can_lehmann_fsm/net430 ),
    .Y(\heichips25_can_lehmann_fsm/_0087_ ),
    .B1(\heichips25_can_lehmann_fsm/_0653_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2376_  (.B1(\heichips25_can_lehmann_fsm/net500 ),
    .Y(\heichips25_can_lehmann_fsm/_0654_ ),
    .A1(\heichips25_can_lehmann_fsm/net983 ),
    .A2(\heichips25_can_lehmann_fsm/net383 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2377_  (.A1(\heichips25_can_lehmann_fsm/_0957_ ),
    .A2(\heichips25_can_lehmann_fsm/net383 ),
    .Y(\heichips25_can_lehmann_fsm/_0088_ ),
    .B1(\heichips25_can_lehmann_fsm/_0654_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2378_  (.B1(\heichips25_can_lehmann_fsm/net495 ),
    .Y(\heichips25_can_lehmann_fsm/_0655_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.const_data[30] ),
    .A2(\heichips25_can_lehmann_fsm/net423 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2379_  (.A1(\heichips25_can_lehmann_fsm/_0957_ ),
    .A2(\heichips25_can_lehmann_fsm/net423 ),
    .Y(\heichips25_can_lehmann_fsm/_0089_ ),
    .B1(\heichips25_can_lehmann_fsm/_0655_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2380_  (.B1(\heichips25_can_lehmann_fsm/net495 ),
    .Y(\heichips25_can_lehmann_fsm/_0656_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.const_data[30] ),
    .A2(\heichips25_can_lehmann_fsm/net382 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2381_  (.A1(\heichips25_can_lehmann_fsm/_0956_ ),
    .A2(\heichips25_can_lehmann_fsm/net382 ),
    .Y(\heichips25_can_lehmann_fsm/_0090_ ),
    .B1(\heichips25_can_lehmann_fsm/_0656_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2382_  (.B1(\heichips25_can_lehmann_fsm/net495 ),
    .Y(\heichips25_can_lehmann_fsm/_0657_ ),
    .A1(\heichips25_can_lehmann_fsm/net912 ),
    .A2(\heichips25_can_lehmann_fsm/net423 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2383_  (.A1(\heichips25_can_lehmann_fsm/_0956_ ),
    .A2(\heichips25_can_lehmann_fsm/net423 ),
    .Y(\heichips25_can_lehmann_fsm/_0091_ ),
    .B1(\heichips25_can_lehmann_fsm/_0657_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2384_  (.B1(\heichips25_can_lehmann_fsm/net481 ),
    .Y(\heichips25_can_lehmann_fsm/_0658_ ),
    .A1(\heichips25_can_lehmann_fsm/net912 ),
    .A2(\heichips25_can_lehmann_fsm/net372 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2385_  (.A1(\heichips25_can_lehmann_fsm/_0955_ ),
    .A2(\heichips25_can_lehmann_fsm/net372 ),
    .Y(\heichips25_can_lehmann_fsm/_0092_ ),
    .B1(\heichips25_can_lehmann_fsm/_0658_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2386_  (.B1(\heichips25_can_lehmann_fsm/net480 ),
    .Y(\heichips25_can_lehmann_fsm/_0659_ ),
    .A1(\heichips25_can_lehmann_fsm/net1068 ),
    .A2(\heichips25_can_lehmann_fsm/net414 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2387_  (.A1(\heichips25_can_lehmann_fsm/_0955_ ),
    .A2(\heichips25_can_lehmann_fsm/net414 ),
    .Y(\heichips25_can_lehmann_fsm/_0093_ ),
    .B1(\heichips25_can_lehmann_fsm/_0659_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2388_  (.B1(\heichips25_can_lehmann_fsm/net480 ),
    .Y(\heichips25_can_lehmann_fsm/_0660_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[34] ),
    .A2(\heichips25_can_lehmann_fsm/net372 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2389_  (.A1(\heichips25_can_lehmann_fsm/_0954_ ),
    .A2(\heichips25_can_lehmann_fsm/net372 ),
    .Y(\heichips25_can_lehmann_fsm/_0094_ ),
    .B1(\heichips25_can_lehmann_fsm/_0660_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2390_  (.B1(\heichips25_can_lehmann_fsm/net480 ),
    .Y(\heichips25_can_lehmann_fsm/_0661_ ),
    .A1(\heichips25_can_lehmann_fsm/net1081 ),
    .A2(\heichips25_can_lehmann_fsm/net399 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2391_  (.A1(\heichips25_can_lehmann_fsm/_0954_ ),
    .A2(\heichips25_can_lehmann_fsm/net399 ),
    .Y(\heichips25_can_lehmann_fsm/_0095_ ),
    .B1(\heichips25_can_lehmann_fsm/_0661_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2392_  (.B1(\heichips25_can_lehmann_fsm/net480 ),
    .Y(\heichips25_can_lehmann_fsm/_0662_ ),
    .A1(\heichips25_can_lehmann_fsm/net1081 ),
    .A2(\heichips25_can_lehmann_fsm/net360 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2393_  (.A1(\heichips25_can_lehmann_fsm/_0953_ ),
    .A2(\heichips25_can_lehmann_fsm/net360 ),
    .Y(\heichips25_can_lehmann_fsm/_0096_ ),
    .B1(\heichips25_can_lehmann_fsm/_0662_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2394_  (.B1(\heichips25_can_lehmann_fsm/net470 ),
    .Y(\heichips25_can_lehmann_fsm/_0663_ ),
    .A1(\heichips25_can_lehmann_fsm/net1066 ),
    .A2(\heichips25_can_lehmann_fsm/net390 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2395_  (.A1(\heichips25_can_lehmann_fsm/_0953_ ),
    .A2(\heichips25_can_lehmann_fsm/net390 ),
    .Y(\heichips25_can_lehmann_fsm/_0097_ ),
    .B1(\heichips25_can_lehmann_fsm/_0663_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2396_  (.B1(\heichips25_can_lehmann_fsm/net470 ),
    .Y(\heichips25_can_lehmann_fsm/_0664_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[39] ),
    .A2(\heichips25_can_lehmann_fsm/net390 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2397_  (.A1(\heichips25_can_lehmann_fsm/_0952_ ),
    .A2(\heichips25_can_lehmann_fsm/net390 ),
    .Y(\heichips25_can_lehmann_fsm/_0098_ ),
    .B1(\heichips25_can_lehmann_fsm/_0664_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2398_  (.B1(\heichips25_can_lehmann_fsm/net470 ),
    .Y(\heichips25_can_lehmann_fsm/_0665_ ),
    .A1(\heichips25_can_lehmann_fsm/net1080 ),
    .A2(\heichips25_can_lehmann_fsm/net355 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2399_  (.A1(\heichips25_can_lehmann_fsm/_0951_ ),
    .A2(\heichips25_can_lehmann_fsm/net355 ),
    .Y(\heichips25_can_lehmann_fsm/_0099_ ),
    .B1(\heichips25_can_lehmann_fsm/_0665_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2400_  (.B1(\heichips25_can_lehmann_fsm/net471 ),
    .Y(\heichips25_can_lehmann_fsm/_0666_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[41] ),
    .A2(\heichips25_can_lehmann_fsm/net402 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2401_  (.A1(\heichips25_can_lehmann_fsm/_0951_ ),
    .A2(\heichips25_can_lehmann_fsm/net390 ),
    .Y(\heichips25_can_lehmann_fsm/_0100_ ),
    .B1(\heichips25_can_lehmann_fsm/_0666_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2402_  (.B1(\heichips25_can_lehmann_fsm/net473 ),
    .Y(\heichips25_can_lehmann_fsm/_0667_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[41] ),
    .A2(\heichips25_can_lehmann_fsm/net364 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2403_  (.A1(\heichips25_can_lehmann_fsm/_0950_ ),
    .A2(\heichips25_can_lehmann_fsm/net364 ),
    .Y(\heichips25_can_lehmann_fsm/_0101_ ),
    .B1(\heichips25_can_lehmann_fsm/_0667_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2404_  (.B1(\heichips25_can_lehmann_fsm/net473 ),
    .Y(\heichips25_can_lehmann_fsm/_0668_ ),
    .A1(\heichips25_can_lehmann_fsm/net1126 ),
    .A2(\heichips25_can_lehmann_fsm/net401 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2405_  (.A1(\heichips25_can_lehmann_fsm/_0950_ ),
    .A2(\heichips25_can_lehmann_fsm/net401 ),
    .Y(\heichips25_can_lehmann_fsm/_0102_ ),
    .B1(\heichips25_can_lehmann_fsm/_0668_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2406_  (.B1(\heichips25_can_lehmann_fsm/net473 ),
    .Y(\heichips25_can_lehmann_fsm/_0669_ ),
    .A1(\heichips25_can_lehmann_fsm/net1055 ),
    .A2(\heichips25_can_lehmann_fsm/net401 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2407_  (.A1(\heichips25_can_lehmann_fsm/_0949_ ),
    .A2(\heichips25_can_lehmann_fsm/net401 ),
    .Y(\heichips25_can_lehmann_fsm/_0103_ ),
    .B1(\heichips25_can_lehmann_fsm/_0669_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2408_  (.B1(\heichips25_can_lehmann_fsm/net493 ),
    .Y(\heichips25_can_lehmann_fsm/_0670_ ),
    .A1(\heichips25_can_lehmann_fsm/net1000 ),
    .A2(\heichips25_can_lehmann_fsm/net405 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2409_  (.A1(\heichips25_can_lehmann_fsm/_0948_ ),
    .A2(\heichips25_can_lehmann_fsm/net405 ),
    .Y(\heichips25_can_lehmann_fsm/_0104_ ),
    .B1(\heichips25_can_lehmann_fsm/_0670_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2410_  (.B1(\heichips25_can_lehmann_fsm/net491 ),
    .Y(\heichips25_can_lehmann_fsm/_0671_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[46] ),
    .A2(\heichips25_can_lehmann_fsm/net421 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2411_  (.A1(\heichips25_can_lehmann_fsm/_0947_ ),
    .A2(\heichips25_can_lehmann_fsm/net421 ),
    .Y(\heichips25_can_lehmann_fsm/_0105_ ),
    .B1(\heichips25_can_lehmann_fsm/_0671_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2412_  (.B1(\heichips25_can_lehmann_fsm/net492 ),
    .Y(\heichips25_can_lehmann_fsm/_0672_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[46] ),
    .A2(\heichips25_can_lehmann_fsm/net380 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2413_  (.A1(\heichips25_can_lehmann_fsm/_0946_ ),
    .A2(\heichips25_can_lehmann_fsm/net380 ),
    .Y(\heichips25_can_lehmann_fsm/_0106_ ),
    .B1(\heichips25_can_lehmann_fsm/_0672_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2414_  (.B1(\heichips25_can_lehmann_fsm/net500 ),
    .Y(\heichips25_can_lehmann_fsm/_0673_ ),
    .A1(\heichips25_can_lehmann_fsm/net879 ),
    .A2(\heichips25_can_lehmann_fsm/net430 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2415_  (.A1(\heichips25_can_lehmann_fsm/_0946_ ),
    .A2(\heichips25_can_lehmann_fsm/net424 ),
    .Y(\heichips25_can_lehmann_fsm/_0107_ ),
    .B1(\heichips25_can_lehmann_fsm/_0673_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2416_  (.B1(\heichips25_can_lehmann_fsm/net499 ),
    .Y(\heichips25_can_lehmann_fsm/_0674_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[49] ),
    .A2(\heichips25_can_lehmann_fsm/net426 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2417_  (.A1(\heichips25_can_lehmann_fsm/_0945_ ),
    .A2(\heichips25_can_lehmann_fsm/net426 ),
    .Y(\heichips25_can_lehmann_fsm/_0108_ ),
    .B1(\heichips25_can_lehmann_fsm/_0674_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2418_  (.B1(\heichips25_can_lehmann_fsm/net497 ),
    .Y(\heichips25_can_lehmann_fsm/_0675_ ),
    .A1(\heichips25_can_lehmann_fsm/net977 ),
    .A2(\heichips25_can_lehmann_fsm/net384 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2419_  (.A1(\heichips25_can_lehmann_fsm/_0944_ ),
    .A2(\heichips25_can_lehmann_fsm/net384 ),
    .Y(\heichips25_can_lehmann_fsm/_0109_ ),
    .B1(\heichips25_can_lehmann_fsm/_0675_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2420_  (.B1(\heichips25_can_lehmann_fsm/net498 ),
    .Y(\heichips25_can_lehmann_fsm/_0676_ ),
    .A1(\heichips25_can_lehmann_fsm/net916 ),
    .A2(\heichips25_can_lehmann_fsm/net427 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2421_  (.A1(\heichips25_can_lehmann_fsm/_0944_ ),
    .A2(\heichips25_can_lehmann_fsm/net427 ),
    .Y(\heichips25_can_lehmann_fsm/_0110_ ),
    .B1(\heichips25_can_lehmann_fsm/_0676_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2422_  (.B1(\heichips25_can_lehmann_fsm/net498 ),
    .Y(\heichips25_can_lehmann_fsm/_0677_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[52] ),
    .A2(\heichips25_can_lehmann_fsm/net427 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2423_  (.A1(\heichips25_can_lehmann_fsm/_0943_ ),
    .A2(\heichips25_can_lehmann_fsm/net427 ),
    .Y(\heichips25_can_lehmann_fsm/_0111_ ),
    .B1(\heichips25_can_lehmann_fsm/_0677_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2424_  (.B1(\heichips25_can_lehmann_fsm/net481 ),
    .Y(\heichips25_can_lehmann_fsm/_0678_ ),
    .A1(\heichips25_can_lehmann_fsm/net1003 ),
    .A2(\heichips25_can_lehmann_fsm/net412 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2425_  (.A1(\heichips25_can_lehmann_fsm/_0942_ ),
    .A2(\heichips25_can_lehmann_fsm/net412 ),
    .Y(\heichips25_can_lehmann_fsm/_0112_ ),
    .B1(\heichips25_can_lehmann_fsm/_0678_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2426_  (.B1(\heichips25_can_lehmann_fsm/net481 ),
    .Y(\heichips25_can_lehmann_fsm/_0679_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[54] ),
    .A2(\heichips25_can_lehmann_fsm/net412 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2427_  (.A1(\heichips25_can_lehmann_fsm/_0941_ ),
    .A2(\heichips25_can_lehmann_fsm/net413 ),
    .Y(\heichips25_can_lehmann_fsm/_0113_ ),
    .B1(\heichips25_can_lehmann_fsm/_0679_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2428_  (.B1(\heichips25_can_lehmann_fsm/net481 ),
    .Y(\heichips25_can_lehmann_fsm/_0680_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[54] ),
    .A2(\heichips25_can_lehmann_fsm/net372 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2429_  (.A1(\heichips25_can_lehmann_fsm/_0940_ ),
    .A2(\heichips25_can_lehmann_fsm/net372 ),
    .Y(\heichips25_can_lehmann_fsm/_0114_ ),
    .B1(\heichips25_can_lehmann_fsm/_0680_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2430_  (.B1(\heichips25_can_lehmann_fsm/net481 ),
    .Y(\heichips25_can_lehmann_fsm/_0681_ ),
    .A1(\heichips25_can_lehmann_fsm/net973 ),
    .A2(\heichips25_can_lehmann_fsm/net412 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2431_  (.A1(\heichips25_can_lehmann_fsm/_0940_ ),
    .A2(\heichips25_can_lehmann_fsm/net412 ),
    .Y(\heichips25_can_lehmann_fsm/_0115_ ),
    .B1(\heichips25_can_lehmann_fsm/_0681_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2432_  (.B1(\heichips25_can_lehmann_fsm/net477 ),
    .Y(\heichips25_can_lehmann_fsm/_0682_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[56] ),
    .A2(\heichips25_can_lehmann_fsm/net370 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2433_  (.A1(\heichips25_can_lehmann_fsm/_0939_ ),
    .A2(\heichips25_can_lehmann_fsm/net370 ),
    .Y(\heichips25_can_lehmann_fsm/_0116_ ),
    .B1(\heichips25_can_lehmann_fsm/_0682_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2434_  (.B1(\heichips25_can_lehmann_fsm/net477 ),
    .Y(\heichips25_can_lehmann_fsm/_0683_ ),
    .A1(\heichips25_can_lehmann_fsm/net989 ),
    .A2(\heichips25_can_lehmann_fsm/net410 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2435_  (.A1(\heichips25_can_lehmann_fsm/_0939_ ),
    .A2(\heichips25_can_lehmann_fsm/net409 ),
    .Y(\heichips25_can_lehmann_fsm/_0117_ ),
    .B1(\heichips25_can_lehmann_fsm/_0683_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2436_  (.B1(\heichips25_can_lehmann_fsm/net477 ),
    .Y(\heichips25_can_lehmann_fsm/_0684_ ),
    .A1(\heichips25_can_lehmann_fsm/net989 ),
    .A2(\heichips25_can_lehmann_fsm/net368 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2437_  (.A1(\heichips25_can_lehmann_fsm/_0938_ ),
    .A2(\heichips25_can_lehmann_fsm/net368 ),
    .Y(\heichips25_can_lehmann_fsm/_0118_ ),
    .B1(\heichips25_can_lehmann_fsm/_0684_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2438_  (.B1(\heichips25_can_lehmann_fsm/net464 ),
    .Y(\heichips25_can_lehmann_fsm/_0685_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[60] ),
    .A2(\heichips25_can_lehmann_fsm/net394 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2439_  (.A1(\heichips25_can_lehmann_fsm/_0938_ ),
    .A2(\heichips25_can_lehmann_fsm/net395 ),
    .Y(\heichips25_can_lehmann_fsm/_0119_ ),
    .B1(\heichips25_can_lehmann_fsm/_0685_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2440_  (.B1(\heichips25_can_lehmann_fsm/net464 ),
    .Y(\heichips25_can_lehmann_fsm/_0686_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[60] ),
    .A2(\heichips25_can_lehmann_fsm/net357 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2441_  (.A1(\heichips25_can_lehmann_fsm/_0937_ ),
    .A2(\heichips25_can_lehmann_fsm/net357 ),
    .Y(\heichips25_can_lehmann_fsm/_0120_ ),
    .B1(\heichips25_can_lehmann_fsm/_0686_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2442_  (.B1(\heichips25_can_lehmann_fsm/net464 ),
    .Y(\heichips25_can_lehmann_fsm/_0687_ ),
    .A1(\heichips25_can_lehmann_fsm/net876 ),
    .A2(\heichips25_can_lehmann_fsm/net394 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2443_  (.A1(\heichips25_can_lehmann_fsm/_0937_ ),
    .A2(\heichips25_can_lehmann_fsm/net394 ),
    .Y(\heichips25_can_lehmann_fsm/_0121_ ),
    .B1(\heichips25_can_lehmann_fsm/_0687_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2444_  (.B1(\heichips25_can_lehmann_fsm/net464 ),
    .Y(\heichips25_can_lehmann_fsm/_0688_ ),
    .A1(\heichips25_can_lehmann_fsm/net876 ),
    .A2(\heichips25_can_lehmann_fsm/net357 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2445_  (.A1(\heichips25_can_lehmann_fsm/_0936_ ),
    .A2(\heichips25_can_lehmann_fsm/net359 ),
    .Y(\heichips25_can_lehmann_fsm/_0122_ ),
    .B1(\heichips25_can_lehmann_fsm/_0688_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2446_  (.B1(\heichips25_can_lehmann_fsm/net468 ),
    .Y(\heichips25_can_lehmann_fsm/_0689_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[64] ),
    .A2(\heichips25_can_lehmann_fsm/net398 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2447_  (.A1(\heichips25_can_lehmann_fsm/_0936_ ),
    .A2(\heichips25_can_lehmann_fsm/net398 ),
    .Y(\heichips25_can_lehmann_fsm/_0123_ ),
    .B1(\heichips25_can_lehmann_fsm/_0689_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2448_  (.B1(\heichips25_can_lehmann_fsm/net468 ),
    .Y(\heichips25_can_lehmann_fsm/_0690_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[64] ),
    .A2(\heichips25_can_lehmann_fsm/net359 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2449_  (.A1(\heichips25_can_lehmann_fsm/_0935_ ),
    .A2(\heichips25_can_lehmann_fsm/net359 ),
    .Y(\heichips25_can_lehmann_fsm/_0124_ ),
    .B1(\heichips25_can_lehmann_fsm/_0690_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2450_  (.B1(\heichips25_can_lehmann_fsm/net468 ),
    .Y(\heichips25_can_lehmann_fsm/_0691_ ),
    .A1(\heichips25_can_lehmann_fsm/net1069 ),
    .A2(\heichips25_can_lehmann_fsm/net398 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2451_  (.A1(\heichips25_can_lehmann_fsm/_0935_ ),
    .A2(\heichips25_can_lehmann_fsm/net398 ),
    .Y(\heichips25_can_lehmann_fsm/_0125_ ),
    .B1(\heichips25_can_lehmann_fsm/_0691_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2452_  (.B1(\heichips25_can_lehmann_fsm/net472 ),
    .Y(\heichips25_can_lehmann_fsm/_0692_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[66] ),
    .A2(\heichips25_can_lehmann_fsm/net365 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2453_  (.A1(\heichips25_can_lehmann_fsm/_0934_ ),
    .A2(\heichips25_can_lehmann_fsm/net365 ),
    .Y(\heichips25_can_lehmann_fsm/_0126_ ),
    .B1(\heichips25_can_lehmann_fsm/_0692_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2454_  (.B1(\heichips25_can_lehmann_fsm/net472 ),
    .Y(\heichips25_can_lehmann_fsm/_0693_ ),
    .A1(\heichips25_can_lehmann_fsm/net1024 ),
    .A2(\heichips25_can_lehmann_fsm/net404 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2455_  (.A1(\heichips25_can_lehmann_fsm/_0934_ ),
    .A2(\heichips25_can_lehmann_fsm/net404 ),
    .Y(\heichips25_can_lehmann_fsm/_0127_ ),
    .B1(\heichips25_can_lehmann_fsm/_0693_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2456_  (.B1(\heichips25_can_lehmann_fsm/net472 ),
    .Y(\heichips25_can_lehmann_fsm/_0694_ ),
    .A1(\heichips25_can_lehmann_fsm/net1024 ),
    .A2(\heichips25_can_lehmann_fsm/net365 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2457_  (.A1(\heichips25_can_lehmann_fsm/_0933_ ),
    .A2(\heichips25_can_lehmann_fsm/net365 ),
    .Y(\heichips25_can_lehmann_fsm/_0128_ ),
    .B1(\heichips25_can_lehmann_fsm/_0694_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2458_  (.B1(\heichips25_can_lehmann_fsm/net493 ),
    .Y(\heichips25_can_lehmann_fsm/_0695_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[70] ),
    .A2(\heichips25_can_lehmann_fsm/net405 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2459_  (.A1(\heichips25_can_lehmann_fsm/_0933_ ),
    .A2(\heichips25_can_lehmann_fsm/net405 ),
    .Y(\heichips25_can_lehmann_fsm/_0129_ ),
    .B1(\heichips25_can_lehmann_fsm/_0695_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2460_  (.B1(\heichips25_can_lehmann_fsm/net492 ),
    .Y(\heichips25_can_lehmann_fsm/_0696_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[70] ),
    .A2(\heichips25_can_lehmann_fsm/net380 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2461_  (.A1(\heichips25_can_lehmann_fsm/_0932_ ),
    .A2(\heichips25_can_lehmann_fsm/net380 ),
    .Y(\heichips25_can_lehmann_fsm/_0130_ ),
    .B1(\heichips25_can_lehmann_fsm/_0696_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2462_  (.B1(\heichips25_can_lehmann_fsm/net499 ),
    .Y(\heichips25_can_lehmann_fsm/_0697_ ),
    .A1(\heichips25_can_lehmann_fsm/net1102 ),
    .A2(\heichips25_can_lehmann_fsm/net429 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2463_  (.A1(\heichips25_can_lehmann_fsm/_0932_ ),
    .A2(\heichips25_can_lehmann_fsm/net422 ),
    .Y(\heichips25_can_lehmann_fsm/_0131_ ),
    .B1(\heichips25_can_lehmann_fsm/_0697_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2464_  (.B1(\heichips25_can_lehmann_fsm/net499 ),
    .Y(\heichips25_can_lehmann_fsm/_0698_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[72] ),
    .A2(\heichips25_can_lehmann_fsm/net386 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2465_  (.A1(\heichips25_can_lehmann_fsm/_0931_ ),
    .A2(\heichips25_can_lehmann_fsm/net386 ),
    .Y(\heichips25_can_lehmann_fsm/_0132_ ),
    .B1(\heichips25_can_lehmann_fsm/_0698_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2466_  (.B1(\heichips25_can_lehmann_fsm/net498 ),
    .Y(\heichips25_can_lehmann_fsm/_0699_ ),
    .A1(\heichips25_can_lehmann_fsm/net903 ),
    .A2(\heichips25_can_lehmann_fsm/net426 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2467_  (.A1(\heichips25_can_lehmann_fsm/_0931_ ),
    .A2(\heichips25_can_lehmann_fsm/net426 ),
    .Y(\heichips25_can_lehmann_fsm/_0133_ ),
    .B1(\heichips25_can_lehmann_fsm/_0699_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2468_  (.B1(\heichips25_can_lehmann_fsm/net498 ),
    .Y(\heichips25_can_lehmann_fsm/_0700_ ),
    .A1(\heichips25_can_lehmann_fsm/net903 ),
    .A2(\heichips25_can_lehmann_fsm/net384 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2469_  (.A1(\heichips25_can_lehmann_fsm/_0930_ ),
    .A2(\heichips25_can_lehmann_fsm/net377 ),
    .Y(\heichips25_can_lehmann_fsm/_0134_ ),
    .B1(\heichips25_can_lehmann_fsm/_0700_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2470_  (.B1(\heichips25_can_lehmann_fsm/net487 ),
    .Y(\heichips25_can_lehmann_fsm/_0701_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[76] ),
    .A2(\heichips25_can_lehmann_fsm/net418 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2471_  (.A1(\heichips25_can_lehmann_fsm/_0930_ ),
    .A2(\heichips25_can_lehmann_fsm/net418 ),
    .Y(\heichips25_can_lehmann_fsm/_0135_ ),
    .B1(\heichips25_can_lehmann_fsm/_0701_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2472_  (.B1(\heichips25_can_lehmann_fsm/net488 ),
    .Y(\heichips25_can_lehmann_fsm/_0702_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[76] ),
    .A2(\heichips25_can_lehmann_fsm/net377 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2473_  (.A1(\heichips25_can_lehmann_fsm/_0929_ ),
    .A2(\heichips25_can_lehmann_fsm/net376 ),
    .Y(\heichips25_can_lehmann_fsm/_0136_ ),
    .B1(\heichips25_can_lehmann_fsm/_0702_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2474_  (.B1(\heichips25_can_lehmann_fsm/net483 ),
    .Y(\heichips25_can_lehmann_fsm/_0703_ ),
    .A1(\heichips25_can_lehmann_fsm/net975 ),
    .A2(\heichips25_can_lehmann_fsm/net415 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2475_  (.A1(\heichips25_can_lehmann_fsm/_0929_ ),
    .A2(\heichips25_can_lehmann_fsm/net415 ),
    .Y(\heichips25_can_lehmann_fsm/_0137_ ),
    .B1(\heichips25_can_lehmann_fsm/_0703_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2476_  (.B1(\heichips25_can_lehmann_fsm/net483 ),
    .Y(\heichips25_can_lehmann_fsm/_0704_ ),
    .A1(\heichips25_can_lehmann_fsm/net975 ),
    .A2(\heichips25_can_lehmann_fsm/net374 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2477_  (.A1(\heichips25_can_lehmann_fsm/_0928_ ),
    .A2(\heichips25_can_lehmann_fsm/net374 ),
    .Y(\heichips25_can_lehmann_fsm/_0138_ ),
    .B1(\heichips25_can_lehmann_fsm/_0704_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2478_  (.B1(\heichips25_can_lehmann_fsm/net483 ),
    .Y(\heichips25_can_lehmann_fsm/_0705_ ),
    .A1(\heichips25_can_lehmann_fsm/net869 ),
    .A2(\heichips25_can_lehmann_fsm/net416 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2479_  (.A1(\heichips25_can_lehmann_fsm/_0928_ ),
    .A2(\heichips25_can_lehmann_fsm/net416 ),
    .Y(\heichips25_can_lehmann_fsm/_0139_ ),
    .B1(\heichips25_can_lehmann_fsm/_0705_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2480_  (.B1(\heichips25_can_lehmann_fsm/net482 ),
    .Y(\heichips25_can_lehmann_fsm/_0706_ ),
    .A1(\heichips25_can_lehmann_fsm/net869 ),
    .A2(\heichips25_can_lehmann_fsm/net370 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2481_  (.A1(\heichips25_can_lehmann_fsm/_0927_ ),
    .A2(\heichips25_can_lehmann_fsm/net370 ),
    .Y(\heichips25_can_lehmann_fsm/_0140_ ),
    .B1(\heichips25_can_lehmann_fsm/_0706_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2482_  (.B1(\heichips25_can_lehmann_fsm/net482 ),
    .Y(\heichips25_can_lehmann_fsm/_0707_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[82] ),
    .A2(\heichips25_can_lehmann_fsm/net409 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2483_  (.A1(\heichips25_can_lehmann_fsm/_0927_ ),
    .A2(\heichips25_can_lehmann_fsm/net409 ),
    .Y(\heichips25_can_lehmann_fsm/_0141_ ),
    .B1(\heichips25_can_lehmann_fsm/_0707_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2484_  (.B1(\heichips25_can_lehmann_fsm/net477 ),
    .Y(\heichips25_can_lehmann_fsm/_0708_ ),
    .A1(\heichips25_can_lehmann_fsm/net1135 ),
    .A2(\heichips25_can_lehmann_fsm/net368 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2485_  (.A1(\heichips25_can_lehmann_fsm/_0926_ ),
    .A2(\heichips25_can_lehmann_fsm/net368 ),
    .Y(\heichips25_can_lehmann_fsm/_0142_ ),
    .B1(\heichips25_can_lehmann_fsm/_0708_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2486_  (.B1(\heichips25_can_lehmann_fsm/net476 ),
    .Y(\heichips25_can_lehmann_fsm/_0709_ ),
    .A1(\heichips25_can_lehmann_fsm/net1070 ),
    .A2(\heichips25_can_lehmann_fsm/net395 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2487_  (.A1(\heichips25_can_lehmann_fsm/_0926_ ),
    .A2(\heichips25_can_lehmann_fsm/net395 ),
    .Y(\heichips25_can_lehmann_fsm/_0143_ ),
    .B1(\heichips25_can_lehmann_fsm/_0709_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2488_  (.B1(\heichips25_can_lehmann_fsm/net464 ),
    .Y(\heichips25_can_lehmann_fsm/_0710_ ),
    .A1(\heichips25_can_lehmann_fsm/net1070 ),
    .A2(\heichips25_can_lehmann_fsm/net358 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2489_  (.A1(\heichips25_can_lehmann_fsm/_0925_ ),
    .A2(\heichips25_can_lehmann_fsm/net357 ),
    .Y(\heichips25_can_lehmann_fsm/_0144_ ),
    .B1(\heichips25_can_lehmann_fsm/_0710_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2490_  (.B1(\heichips25_can_lehmann_fsm/net464 ),
    .Y(\heichips25_can_lehmann_fsm/_0711_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[86] ),
    .A2(\heichips25_can_lehmann_fsm/net394 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2491_  (.A1(\heichips25_can_lehmann_fsm/_0925_ ),
    .A2(\heichips25_can_lehmann_fsm/net394 ),
    .Y(\heichips25_can_lehmann_fsm/_0145_ ),
    .B1(\heichips25_can_lehmann_fsm/_0711_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2492_  (.B1(\heichips25_can_lehmann_fsm/net466 ),
    .Y(\heichips25_can_lehmann_fsm/_0712_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[86] ),
    .A2(\heichips25_can_lehmann_fsm/net356 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2493_  (.A1(\heichips25_can_lehmann_fsm/_0924_ ),
    .A2(\heichips25_can_lehmann_fsm/net356 ),
    .Y(\heichips25_can_lehmann_fsm/_0146_ ),
    .B1(\heichips25_can_lehmann_fsm/_0712_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2494_  (.B1(\heichips25_can_lehmann_fsm/net467 ),
    .Y(\heichips25_can_lehmann_fsm/_0713_ ),
    .A1(\heichips25_can_lehmann_fsm/net962 ),
    .A2(\heichips25_can_lehmann_fsm/net390 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2495_  (.A1(\heichips25_can_lehmann_fsm/_0924_ ),
    .A2(\heichips25_can_lehmann_fsm/net390 ),
    .Y(\heichips25_can_lehmann_fsm/_0147_ ),
    .B1(\heichips25_can_lehmann_fsm/_0713_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2496_  (.B1(\heichips25_can_lehmann_fsm/net467 ),
    .Y(\heichips25_can_lehmann_fsm/_0714_ ),
    .A1(\heichips25_can_lehmann_fsm/net962 ),
    .A2(\heichips25_can_lehmann_fsm/net355 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2497_  (.A1(\heichips25_can_lehmann_fsm/_0923_ ),
    .A2(\heichips25_can_lehmann_fsm/net355 ),
    .Y(\heichips25_can_lehmann_fsm/_0148_ ),
    .B1(\heichips25_can_lehmann_fsm/_0714_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2498_  (.B1(\heichips25_can_lehmann_fsm/net467 ),
    .Y(\heichips25_can_lehmann_fsm/_0715_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[90] ),
    .A2(\heichips25_can_lehmann_fsm/net391 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2499_  (.A1(\heichips25_can_lehmann_fsm/_0923_ ),
    .A2(\heichips25_can_lehmann_fsm/net391 ),
    .Y(\heichips25_can_lehmann_fsm/_0149_ ),
    .B1(\heichips25_can_lehmann_fsm/_0715_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2500_  (.B1(\heichips25_can_lehmann_fsm/net469 ),
    .Y(\heichips25_can_lehmann_fsm/_0716_ ),
    .A1(\heichips25_can_lehmann_fsm/net1054 ),
    .A2(\heichips25_can_lehmann_fsm/net359 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2501_  (.A1(\heichips25_can_lehmann_fsm/_0922_ ),
    .A2(\heichips25_can_lehmann_fsm/net359 ),
    .Y(\heichips25_can_lehmann_fsm/_0150_ ),
    .B1(\heichips25_can_lehmann_fsm/_0716_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2502_  (.B1(\heichips25_can_lehmann_fsm/net493 ),
    .Y(\heichips25_can_lehmann_fsm/_0717_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[92] ),
    .A2(\heichips25_can_lehmann_fsm/net405 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2503_  (.A1(\heichips25_can_lehmann_fsm/_0922_ ),
    .A2(\heichips25_can_lehmann_fsm/net407 ),
    .Y(\heichips25_can_lehmann_fsm/_0151_ ),
    .B1(\heichips25_can_lehmann_fsm/_0717_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2504_  (.B1(\heichips25_can_lehmann_fsm/net493 ),
    .Y(\heichips25_can_lehmann_fsm/_0718_ ),
    .A1(\heichips25_can_lehmann_fsm/net1092 ),
    .A2(\heichips25_can_lehmann_fsm/net366 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2505_  (.A1(\heichips25_can_lehmann_fsm/_0921_ ),
    .A2(\heichips25_can_lehmann_fsm/net366 ),
    .Y(\heichips25_can_lehmann_fsm/_0152_ ),
    .B1(\heichips25_can_lehmann_fsm/_0718_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2506_  (.B1(\heichips25_can_lehmann_fsm/net491 ),
    .Y(\heichips25_can_lehmann_fsm/_0719_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[94] ),
    .A2(\heichips25_can_lehmann_fsm/net421 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2507_  (.A1(\heichips25_can_lehmann_fsm/_0921_ ),
    .A2(\heichips25_can_lehmann_fsm/net421 ),
    .Y(\heichips25_can_lehmann_fsm/_0153_ ),
    .B1(\heichips25_can_lehmann_fsm/_0719_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2508_  (.B1(\heichips25_can_lehmann_fsm/net492 ),
    .Y(\heichips25_can_lehmann_fsm/_0720_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[94] ),
    .A2(\heichips25_can_lehmann_fsm/net380 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2509_  (.A1(\heichips25_can_lehmann_fsm/_0920_ ),
    .A2(\heichips25_can_lehmann_fsm/net381 ),
    .Y(\heichips25_can_lehmann_fsm/_0154_ ),
    .B1(\heichips25_can_lehmann_fsm/_0720_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2510_  (.B1(\heichips25_can_lehmann_fsm/net499 ),
    .Y(\heichips25_can_lehmann_fsm/_0721_ ),
    .A1(\heichips25_can_lehmann_fsm/net936 ),
    .A2(\heichips25_can_lehmann_fsm/net422 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2511_  (.A1(\heichips25_can_lehmann_fsm/_0920_ ),
    .A2(\heichips25_can_lehmann_fsm/net422 ),
    .Y(\heichips25_can_lehmann_fsm/_0155_ ),
    .B1(\heichips25_can_lehmann_fsm/_0721_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2512_  (.B1(\heichips25_can_lehmann_fsm/net499 ),
    .Y(\heichips25_can_lehmann_fsm/_0722_ ),
    .A1(\heichips25_can_lehmann_fsm/net936 ),
    .A2(\heichips25_can_lehmann_fsm/net386 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2513_  (.A1(\heichips25_can_lehmann_fsm/_0919_ ),
    .A2(\heichips25_can_lehmann_fsm/net386 ),
    .Y(\heichips25_can_lehmann_fsm/_0156_ ),
    .B1(\heichips25_can_lehmann_fsm/_0722_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2514_  (.B1(\heichips25_can_lehmann_fsm/net499 ),
    .Y(\heichips25_can_lehmann_fsm/_0723_ ),
    .A1(\heichips25_can_lehmann_fsm/net950 ),
    .A2(\heichips25_can_lehmann_fsm/net426 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2515_  (.A1(\heichips25_can_lehmann_fsm/_0919_ ),
    .A2(\heichips25_can_lehmann_fsm/net426 ),
    .Y(\heichips25_can_lehmann_fsm/_0157_ ),
    .B1(\heichips25_can_lehmann_fsm/_0723_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2516_  (.B1(\heichips25_can_lehmann_fsm/net485 ),
    .Y(\heichips25_can_lehmann_fsm/_0724_ ),
    .A1(\heichips25_can_lehmann_fsm/net950 ),
    .A2(\heichips25_can_lehmann_fsm/net378 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2517_  (.A1(\heichips25_can_lehmann_fsm/_0918_ ),
    .A2(\heichips25_can_lehmann_fsm/net378 ),
    .Y(\heichips25_can_lehmann_fsm/_0158_ ),
    .B1(\heichips25_can_lehmann_fsm/_0724_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2518_  (.B1(\heichips25_can_lehmann_fsm/net485 ),
    .Y(\heichips25_can_lehmann_fsm/_0725_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[100] ),
    .A2(\heichips25_can_lehmann_fsm/net417 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2519_  (.A1(\heichips25_can_lehmann_fsm/_0918_ ),
    .A2(\heichips25_can_lehmann_fsm/net417 ),
    .Y(\heichips25_can_lehmann_fsm/_0159_ ),
    .B1(\heichips25_can_lehmann_fsm/_0725_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2520_  (.B1(\heichips25_can_lehmann_fsm/net487 ),
    .Y(\heichips25_can_lehmann_fsm/_0726_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[100] ),
    .A2(\heichips25_can_lehmann_fsm/net378 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2521_  (.A1(\heichips25_can_lehmann_fsm/_0917_ ),
    .A2(\heichips25_can_lehmann_fsm/net376 ),
    .Y(\heichips25_can_lehmann_fsm/_0160_ ),
    .B1(\heichips25_can_lehmann_fsm/_0726_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2522_  (.B1(\heichips25_can_lehmann_fsm/net483 ),
    .Y(\heichips25_can_lehmann_fsm/_0727_ ),
    .A1(\heichips25_can_lehmann_fsm/net1079 ),
    .A2(\heichips25_can_lehmann_fsm/net415 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2523_  (.A1(\heichips25_can_lehmann_fsm/_0917_ ),
    .A2(\heichips25_can_lehmann_fsm/net415 ),
    .Y(\heichips25_can_lehmann_fsm/_0161_ ),
    .B1(\heichips25_can_lehmann_fsm/_0727_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2524_  (.B1(\heichips25_can_lehmann_fsm/net483 ),
    .Y(\heichips25_can_lehmann_fsm/_0728_ ),
    .A1(\heichips25_can_lehmann_fsm/net1079 ),
    .A2(\heichips25_can_lehmann_fsm/net375 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2525_  (.A1(\heichips25_can_lehmann_fsm/_0916_ ),
    .A2(\heichips25_can_lehmann_fsm/net375 ),
    .Y(\heichips25_can_lehmann_fsm/_0162_ ),
    .B1(\heichips25_can_lehmann_fsm/_0728_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2526_  (.B1(\heichips25_can_lehmann_fsm/net483 ),
    .Y(\heichips25_can_lehmann_fsm/_0729_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[104] ),
    .A2(\heichips25_can_lehmann_fsm/net415 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2527_  (.A1(\heichips25_can_lehmann_fsm/_0916_ ),
    .A2(\heichips25_can_lehmann_fsm/net415 ),
    .Y(\heichips25_can_lehmann_fsm/_0163_ ),
    .B1(\heichips25_can_lehmann_fsm/_0729_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2528_  (.B1(\heichips25_can_lehmann_fsm/net477 ),
    .Y(\heichips25_can_lehmann_fsm/_0730_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[104] ),
    .A2(\heichips25_can_lehmann_fsm/net370 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2529_  (.A1(\heichips25_can_lehmann_fsm/_0915_ ),
    .A2(\heichips25_can_lehmann_fsm/net370 ),
    .Y(\heichips25_can_lehmann_fsm/_0164_ ),
    .B1(\heichips25_can_lehmann_fsm/_0730_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2530_  (.B1(\heichips25_can_lehmann_fsm/net478 ),
    .Y(\heichips25_can_lehmann_fsm/_0731_ ),
    .A1(\heichips25_can_lehmann_fsm/net1005 ),
    .A2(\heichips25_can_lehmann_fsm/net410 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2531_  (.A1(\heichips25_can_lehmann_fsm/_0915_ ),
    .A2(\heichips25_can_lehmann_fsm/net409 ),
    .Y(\heichips25_can_lehmann_fsm/_0165_ ),
    .B1(\heichips25_can_lehmann_fsm/_0731_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2532_  (.B1(\heichips25_can_lehmann_fsm/net477 ),
    .Y(\heichips25_can_lehmann_fsm/_0732_ ),
    .A1(\heichips25_can_lehmann_fsm/net1005 ),
    .A2(\heichips25_can_lehmann_fsm/net368 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2533_  (.A1(\heichips25_can_lehmann_fsm/_0914_ ),
    .A2(\heichips25_can_lehmann_fsm/net368 ),
    .Y(\heichips25_can_lehmann_fsm/_0166_ ),
    .B1(\heichips25_can_lehmann_fsm/_0732_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2534_  (.B1(\heichips25_can_lehmann_fsm/net476 ),
    .Y(\heichips25_can_lehmann_fsm/_0733_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[108] ),
    .A2(\heichips25_can_lehmann_fsm/net395 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2535_  (.A1(\heichips25_can_lehmann_fsm/_0914_ ),
    .A2(\heichips25_can_lehmann_fsm/net395 ),
    .Y(\heichips25_can_lehmann_fsm/_0167_ ),
    .B1(\heichips25_can_lehmann_fsm/_0733_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2536_  (.B1(\heichips25_can_lehmann_fsm/net476 ),
    .Y(\heichips25_can_lehmann_fsm/_0734_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[108] ),
    .A2(\heichips25_can_lehmann_fsm/net358 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2537_  (.A1(\heichips25_can_lehmann_fsm/_0913_ ),
    .A2(\heichips25_can_lehmann_fsm/net357 ),
    .Y(\heichips25_can_lehmann_fsm/_0168_ ),
    .B1(\heichips25_can_lehmann_fsm/_0734_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2538_  (.B1(\heichips25_can_lehmann_fsm/net466 ),
    .Y(\heichips25_can_lehmann_fsm/_0735_ ),
    .A1(\heichips25_can_lehmann_fsm/net969 ),
    .A2(\heichips25_can_lehmann_fsm/net393 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2539_  (.A1(\heichips25_can_lehmann_fsm/_0913_ ),
    .A2(\heichips25_can_lehmann_fsm/net393 ),
    .Y(\heichips25_can_lehmann_fsm/_0169_ ),
    .B1(\heichips25_can_lehmann_fsm/_0735_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2540_  (.B1(\heichips25_can_lehmann_fsm/net466 ),
    .Y(\heichips25_can_lehmann_fsm/_0736_ ),
    .A1(\heichips25_can_lehmann_fsm/net969 ),
    .A2(\heichips25_can_lehmann_fsm/net356 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2541_  (.A1(\heichips25_can_lehmann_fsm/_0912_ ),
    .A2(\heichips25_can_lehmann_fsm/net356 ),
    .Y(\heichips25_can_lehmann_fsm/_0170_ ),
    .B1(\heichips25_can_lehmann_fsm/_0736_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2542_  (.B1(\heichips25_can_lehmann_fsm/net467 ),
    .Y(\heichips25_can_lehmann_fsm/_0737_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[112] ),
    .A2(\heichips25_can_lehmann_fsm/net392 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2543_  (.A1(\heichips25_can_lehmann_fsm/_0912_ ),
    .A2(\heichips25_can_lehmann_fsm/net392 ),
    .Y(\heichips25_can_lehmann_fsm/_0171_ ),
    .B1(\heichips25_can_lehmann_fsm/_0737_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2544_  (.B1(\heichips25_can_lehmann_fsm/net467 ),
    .Y(\heichips25_can_lehmann_fsm/_0738_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[112] ),
    .A2(\heichips25_can_lehmann_fsm/net355 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2545_  (.A1(\heichips25_can_lehmann_fsm/_0911_ ),
    .A2(\heichips25_can_lehmann_fsm/net355 ),
    .Y(\heichips25_can_lehmann_fsm/_0172_ ),
    .B1(\heichips25_can_lehmann_fsm/_0738_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2546_  (.B1(\heichips25_can_lehmann_fsm/net467 ),
    .Y(\heichips25_can_lehmann_fsm/_0739_ ),
    .A1(\heichips25_can_lehmann_fsm/net1037 ),
    .A2(\heichips25_can_lehmann_fsm/net392 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2547_  (.A1(\heichips25_can_lehmann_fsm/_0911_ ),
    .A2(\heichips25_can_lehmann_fsm/net392 ),
    .Y(\heichips25_can_lehmann_fsm/_0173_ ),
    .B1(\heichips25_can_lehmann_fsm/_0739_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2548_  (.B1(\heichips25_can_lehmann_fsm/net473 ),
    .Y(\heichips25_can_lehmann_fsm/_0740_ ),
    .A1(\heichips25_can_lehmann_fsm/net1037 ),
    .A2(\heichips25_can_lehmann_fsm/net364 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2549_  (.A1(\heichips25_can_lehmann_fsm/_0910_ ),
    .A2(\heichips25_can_lehmann_fsm/net364 ),
    .Y(\heichips25_can_lehmann_fsm/_0174_ ),
    .B1(\heichips25_can_lehmann_fsm/_0740_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2550_  (.B1(\heichips25_can_lehmann_fsm/net473 ),
    .Y(\heichips25_can_lehmann_fsm/_0741_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[116] ),
    .A2(\heichips25_can_lehmann_fsm/net402 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2551_  (.A1(\heichips25_can_lehmann_fsm/_0910_ ),
    .A2(\heichips25_can_lehmann_fsm/net402 ),
    .Y(\heichips25_can_lehmann_fsm/_0175_ ),
    .B1(\heichips25_can_lehmann_fsm/_0741_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2552_  (.B1(\heichips25_can_lehmann_fsm/net472 ),
    .Y(\heichips25_can_lehmann_fsm/_0742_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[116] ),
    .A2(\heichips25_can_lehmann_fsm/net365 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2553_  (.A1(\heichips25_can_lehmann_fsm/_0909_ ),
    .A2(\heichips25_can_lehmann_fsm/net367 ),
    .Y(\heichips25_can_lehmann_fsm/_0176_ ),
    .B1(\heichips25_can_lehmann_fsm/_0742_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2554_  (.B1(\heichips25_can_lehmann_fsm/net494 ),
    .Y(\heichips25_can_lehmann_fsm/_0743_ ),
    .A1(\heichips25_can_lehmann_fsm/net1082 ),
    .A2(\heichips25_can_lehmann_fsm/net407 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2555_  (.A1(\heichips25_can_lehmann_fsm/_0909_ ),
    .A2(\heichips25_can_lehmann_fsm/net407 ),
    .Y(\heichips25_can_lehmann_fsm/_0177_ ),
    .B1(\heichips25_can_lehmann_fsm/_0743_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2556_  (.B1(\heichips25_can_lehmann_fsm/net495 ),
    .Y(\heichips25_can_lehmann_fsm/_0744_ ),
    .A1(\heichips25_can_lehmann_fsm/net1082 ),
    .A2(\heichips25_can_lehmann_fsm/net382 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2557_  (.A1(\heichips25_can_lehmann_fsm/_0908_ ),
    .A2(\heichips25_can_lehmann_fsm/net382 ),
    .Y(\heichips25_can_lehmann_fsm/_0178_ ),
    .B1(\heichips25_can_lehmann_fsm/_0744_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2558_  (.B1(\heichips25_can_lehmann_fsm/net500 ),
    .Y(\heichips25_can_lehmann_fsm/_0745_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[120] ),
    .A2(\heichips25_can_lehmann_fsm/net430 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2559_  (.A1(\heichips25_can_lehmann_fsm/_0908_ ),
    .A2(\heichips25_can_lehmann_fsm/net430 ),
    .Y(\heichips25_can_lehmann_fsm/_0179_ ),
    .B1(\heichips25_can_lehmann_fsm/_0745_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2560_  (.B1(\heichips25_can_lehmann_fsm/net497 ),
    .Y(\heichips25_can_lehmann_fsm/_0746_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[120] ),
    .A2(\heichips25_can_lehmann_fsm/net386 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2561_  (.A1(\heichips25_can_lehmann_fsm/_0907_ ),
    .A2(\heichips25_can_lehmann_fsm/net386 ),
    .Y(\heichips25_can_lehmann_fsm/_0180_ ),
    .B1(\heichips25_can_lehmann_fsm/_0746_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2562_  (.B1(\heichips25_can_lehmann_fsm/net497 ),
    .Y(\heichips25_can_lehmann_fsm/_0747_ ),
    .A1(\heichips25_can_lehmann_fsm/net1040 ),
    .A2(\heichips25_can_lehmann_fsm/net427 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2563_  (.A1(\heichips25_can_lehmann_fsm/_0907_ ),
    .A2(\heichips25_can_lehmann_fsm/net427 ),
    .Y(\heichips25_can_lehmann_fsm/_0181_ ),
    .B1(\heichips25_can_lehmann_fsm/_0747_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2564_  (.B1(\heichips25_can_lehmann_fsm/net488 ),
    .Y(\heichips25_can_lehmann_fsm/_0748_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[122] ),
    .A2(\heichips25_can_lehmann_fsm/net377 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2565_  (.A1(\heichips25_can_lehmann_fsm/_0906_ ),
    .A2(\heichips25_can_lehmann_fsm/net377 ),
    .Y(\heichips25_can_lehmann_fsm/_0182_ ),
    .B1(\heichips25_can_lehmann_fsm/_0748_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2566_  (.B1(\heichips25_can_lehmann_fsm/net488 ),
    .Y(\heichips25_can_lehmann_fsm/_0749_ ),
    .A1(\heichips25_can_lehmann_fsm/net1109 ),
    .A2(\heichips25_can_lehmann_fsm/net418 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2567_  (.A1(\heichips25_can_lehmann_fsm/_0906_ ),
    .A2(\heichips25_can_lehmann_fsm/net418 ),
    .Y(\heichips25_can_lehmann_fsm/_0183_ ),
    .B1(\heichips25_can_lehmann_fsm/_0749_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2568_  (.B1(\heichips25_can_lehmann_fsm/net487 ),
    .Y(\heichips25_can_lehmann_fsm/_0750_ ),
    .A1(\heichips25_can_lehmann_fsm/net1109 ),
    .A2(\heichips25_can_lehmann_fsm/net376 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2569_  (.A1(\heichips25_can_lehmann_fsm/_0905_ ),
    .A2(\heichips25_can_lehmann_fsm/net376 ),
    .Y(\heichips25_can_lehmann_fsm/_0184_ ),
    .B1(\heichips25_can_lehmann_fsm/_0750_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2570_  (.B1(\heichips25_can_lehmann_fsm/net487 ),
    .Y(\heichips25_can_lehmann_fsm/_0751_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[126] ),
    .A2(\heichips25_can_lehmann_fsm/net418 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2571_  (.A1(\heichips25_can_lehmann_fsm/_0905_ ),
    .A2(\heichips25_can_lehmann_fsm/net418 ),
    .Y(\heichips25_can_lehmann_fsm/_0185_ ),
    .B1(\heichips25_can_lehmann_fsm/_0751_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2572_  (.B1(\heichips25_can_lehmann_fsm/net482 ),
    .Y(\heichips25_can_lehmann_fsm/_0752_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[126] ),
    .A2(\heichips25_can_lehmann_fsm/net374 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2573_  (.A1(\heichips25_can_lehmann_fsm/_0904_ ),
    .A2(\heichips25_can_lehmann_fsm/net374 ),
    .Y(\heichips25_can_lehmann_fsm/_0186_ ),
    .B1(\heichips25_can_lehmann_fsm/_0752_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2574_  (.B1(\heichips25_can_lehmann_fsm/net482 ),
    .Y(\heichips25_can_lehmann_fsm/_0753_ ),
    .A1(\heichips25_can_lehmann_fsm/net1038 ),
    .A2(\heichips25_can_lehmann_fsm/net409 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2575_  (.A1(\heichips25_can_lehmann_fsm/_0904_ ),
    .A2(\heichips25_can_lehmann_fsm/net409 ),
    .Y(\heichips25_can_lehmann_fsm/_0187_ ),
    .B1(\heichips25_can_lehmann_fsm/_0753_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2576_  (.B1(\heichips25_can_lehmann_fsm/net482 ),
    .Y(\heichips25_can_lehmann_fsm/_0754_ ),
    .A1(\heichips25_can_lehmann_fsm/net1038 ),
    .A2(\heichips25_can_lehmann_fsm/net370 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2577_  (.A1(\heichips25_can_lehmann_fsm/_0903_ ),
    .A2(\heichips25_can_lehmann_fsm/net370 ),
    .Y(\heichips25_can_lehmann_fsm/_0188_ ),
    .B1(\heichips25_can_lehmann_fsm/_0754_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2578_  (.B1(\heichips25_can_lehmann_fsm/net478 ),
    .Y(\heichips25_can_lehmann_fsm/_0755_ ),
    .A1(\heichips25_can_lehmann_fsm/net1091 ),
    .A2(\heichips25_can_lehmann_fsm/net411 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2579_  (.A1(\heichips25_can_lehmann_fsm/_0903_ ),
    .A2(\heichips25_can_lehmann_fsm/net411 ),
    .Y(\heichips25_can_lehmann_fsm/_0189_ ),
    .B1(\heichips25_can_lehmann_fsm/_0755_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2580_  (.B1(\heichips25_can_lehmann_fsm/net478 ),
    .Y(\heichips25_can_lehmann_fsm/_0756_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[130] ),
    .A2(\heichips25_can_lehmann_fsm/net369 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2581_  (.A1(\heichips25_can_lehmann_fsm/_0902_ ),
    .A2(\heichips25_can_lehmann_fsm/net369 ),
    .Y(\heichips25_can_lehmann_fsm/_0190_ ),
    .B1(\heichips25_can_lehmann_fsm/_0756_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2582_  (.B1(\heichips25_can_lehmann_fsm/net476 ),
    .Y(\heichips25_can_lehmann_fsm/_0757_ ),
    .A1(\heichips25_can_lehmann_fsm/net902 ),
    .A2(\heichips25_can_lehmann_fsm/net410 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2583_  (.A1(\heichips25_can_lehmann_fsm/_0902_ ),
    .A2(\heichips25_can_lehmann_fsm/net410 ),
    .Y(\heichips25_can_lehmann_fsm/_0191_ ),
    .B1(\heichips25_can_lehmann_fsm/_0757_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2584_  (.B1(\heichips25_can_lehmann_fsm/net476 ),
    .Y(\heichips25_can_lehmann_fsm/_0758_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[132] ),
    .A2(\heichips25_can_lehmann_fsm/net358 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2585_  (.A1(\heichips25_can_lehmann_fsm/_0901_ ),
    .A2(\heichips25_can_lehmann_fsm/net358 ),
    .Y(\heichips25_can_lehmann_fsm/_0192_ ),
    .B1(\heichips25_can_lehmann_fsm/_0758_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2586_  (.B1(\heichips25_can_lehmann_fsm/net476 ),
    .Y(\heichips25_can_lehmann_fsm/_0759_ ),
    .A1(\heichips25_can_lehmann_fsm/net921 ),
    .A2(\heichips25_can_lehmann_fsm/net396 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2587_  (.A1(\heichips25_can_lehmann_fsm/_0901_ ),
    .A2(\heichips25_can_lehmann_fsm/net396 ),
    .Y(\heichips25_can_lehmann_fsm/_0193_ ),
    .B1(\heichips25_can_lehmann_fsm/_0759_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2588_  (.B1(\heichips25_can_lehmann_fsm/net476 ),
    .Y(\heichips25_can_lehmann_fsm/_0760_ ),
    .A1(\heichips25_can_lehmann_fsm/net921 ),
    .A2(\heichips25_can_lehmann_fsm/net358 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2589_  (.A1(\heichips25_can_lehmann_fsm/_0900_ ),
    .A2(\heichips25_can_lehmann_fsm/net360 ),
    .Y(\heichips25_can_lehmann_fsm/_0194_ ),
    .B1(\heichips25_can_lehmann_fsm/_0760_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2590_  (.B1(\heichips25_can_lehmann_fsm/net480 ),
    .Y(\heichips25_can_lehmann_fsm/_0761_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[136] ),
    .A2(\heichips25_can_lehmann_fsm/net399 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2591_  (.A1(\heichips25_can_lehmann_fsm/_0900_ ),
    .A2(\heichips25_can_lehmann_fsm/net399 ),
    .Y(\heichips25_can_lehmann_fsm/_0195_ ),
    .B1(\heichips25_can_lehmann_fsm/_0761_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2592_  (.B1(\heichips25_can_lehmann_fsm/net468 ),
    .Y(\heichips25_can_lehmann_fsm/_0762_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[136] ),
    .A2(\heichips25_can_lehmann_fsm/net360 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2593_  (.A1(\heichips25_can_lehmann_fsm/_0899_ ),
    .A2(\heichips25_can_lehmann_fsm/net360 ),
    .Y(\heichips25_can_lehmann_fsm/_0196_ ),
    .B1(\heichips25_can_lehmann_fsm/_0762_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2594_  (.B1(\heichips25_can_lehmann_fsm/net480 ),
    .Y(\heichips25_can_lehmann_fsm/_0763_ ),
    .A1(\heichips25_can_lehmann_fsm/net972 ),
    .A2(\heichips25_can_lehmann_fsm/net399 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2595_  (.A1(\heichips25_can_lehmann_fsm/_0899_ ),
    .A2(\heichips25_can_lehmann_fsm/net400 ),
    .Y(\heichips25_can_lehmann_fsm/_0197_ ),
    .B1(\heichips25_can_lehmann_fsm/_0763_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2596_  (.B1(\heichips25_can_lehmann_fsm/net480 ),
    .Y(\heichips25_can_lehmann_fsm/_0764_ ),
    .A1(\heichips25_can_lehmann_fsm/net972 ),
    .A2(\heichips25_can_lehmann_fsm/net360 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2597_  (.A1(\heichips25_can_lehmann_fsm/_0898_ ),
    .A2(\heichips25_can_lehmann_fsm/net366 ),
    .Y(\heichips25_can_lehmann_fsm/_0198_ ),
    .B1(\heichips25_can_lehmann_fsm/_0764_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2598_  (.B1(\heichips25_can_lehmann_fsm/net493 ),
    .Y(\heichips25_can_lehmann_fsm/_0765_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[140] ),
    .A2(\heichips25_can_lehmann_fsm/net407 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2599_  (.A1(\heichips25_can_lehmann_fsm/_0898_ ),
    .A2(\heichips25_can_lehmann_fsm/net407 ),
    .Y(\heichips25_can_lehmann_fsm/_0199_ ),
    .B1(\heichips25_can_lehmann_fsm/_0765_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2600_  (.B1(\heichips25_can_lehmann_fsm/net493 ),
    .Y(\heichips25_can_lehmann_fsm/_0766_ ),
    .A1(\heichips25_can_lehmann_fsm/net959 ),
    .A2(\heichips25_can_lehmann_fsm/net366 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2601_  (.A1(\heichips25_can_lehmann_fsm/_0897_ ),
    .A2(\heichips25_can_lehmann_fsm/net366 ),
    .Y(\heichips25_can_lehmann_fsm/_0200_ ),
    .B1(\heichips25_can_lehmann_fsm/_0766_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2602_  (.B1(\heichips25_can_lehmann_fsm/net493 ),
    .Y(\heichips25_can_lehmann_fsm/_0767_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[142] ),
    .A2(\heichips25_can_lehmann_fsm/net422 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2603_  (.A1(\heichips25_can_lehmann_fsm/_0897_ ),
    .A2(\heichips25_can_lehmann_fsm/net422 ),
    .Y(\heichips25_can_lehmann_fsm/_0201_ ),
    .B1(\heichips25_can_lehmann_fsm/_0767_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2604_  (.B1(\heichips25_can_lehmann_fsm/net491 ),
    .Y(\heichips25_can_lehmann_fsm/_0768_ ),
    .A1(\heichips25_can_lehmann_fsm/net930 ),
    .A2(\heichips25_can_lehmann_fsm/net380 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2605_  (.A1(\heichips25_can_lehmann_fsm/_0896_ ),
    .A2(\heichips25_can_lehmann_fsm/net380 ),
    .Y(\heichips25_can_lehmann_fsm/_0202_ ),
    .B1(\heichips25_can_lehmann_fsm/_0768_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2606_  (.B1(\heichips25_can_lehmann_fsm/net491 ),
    .Y(\heichips25_can_lehmann_fsm/_0769_ ),
    .A1(\heichips25_can_lehmann_fsm/net897 ),
    .A2(\heichips25_can_lehmann_fsm/net422 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2607_  (.A1(\heichips25_can_lehmann_fsm/_0896_ ),
    .A2(\heichips25_can_lehmann_fsm/net422 ),
    .Y(\heichips25_can_lehmann_fsm/_0203_ ),
    .B1(\heichips25_can_lehmann_fsm/_0769_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2608_  (.B1(\heichips25_can_lehmann_fsm/net499 ),
    .Y(\heichips25_can_lehmann_fsm/_0770_ ),
    .A1(\heichips25_can_lehmann_fsm/net897 ),
    .A2(\heichips25_can_lehmann_fsm/net381 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2609_  (.A1(\heichips25_can_lehmann_fsm/_0895_ ),
    .A2(\heichips25_can_lehmann_fsm/net381 ),
    .Y(\heichips25_can_lehmann_fsm/_0204_ ),
    .B1(\heichips25_can_lehmann_fsm/_0770_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2610_  (.B1(\heichips25_can_lehmann_fsm/net485 ),
    .Y(\heichips25_can_lehmann_fsm/_0771_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[146] ),
    .A2(\heichips25_can_lehmann_fsm/net413 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2611_  (.A1(\heichips25_can_lehmann_fsm/_0895_ ),
    .A2(\heichips25_can_lehmann_fsm/net425 ),
    .Y(\heichips25_can_lehmann_fsm/_0205_ ),
    .B1(\heichips25_can_lehmann_fsm/_0771_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2612_  (.B1(\heichips25_can_lehmann_fsm/net485 ),
    .Y(\heichips25_can_lehmann_fsm/_0772_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[146] ),
    .A2(\heichips25_can_lehmann_fsm/net372 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2613_  (.A1(\heichips25_can_lehmann_fsm/_0894_ ),
    .A2(\heichips25_can_lehmann_fsm/net372 ),
    .Y(\heichips25_can_lehmann_fsm/_0206_ ),
    .B1(\heichips25_can_lehmann_fsm/_0772_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2614_  (.B1(\heichips25_can_lehmann_fsm/net486 ),
    .Y(\heichips25_can_lehmann_fsm/_0773_ ),
    .A1(\heichips25_can_lehmann_fsm/net1030 ),
    .A2(\heichips25_can_lehmann_fsm/net413 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2615_  (.A1(\heichips25_can_lehmann_fsm/_0894_ ),
    .A2(\heichips25_can_lehmann_fsm/net413 ),
    .Y(\heichips25_can_lehmann_fsm/_0207_ ),
    .B1(\heichips25_can_lehmann_fsm/_0773_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2616_  (.B1(\heichips25_can_lehmann_fsm/net486 ),
    .Y(\heichips25_can_lehmann_fsm/_0774_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[148] ),
    .A2(\heichips25_can_lehmann_fsm/net373 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2617_  (.A1(\heichips25_can_lehmann_fsm/_0893_ ),
    .A2(\heichips25_can_lehmann_fsm/net373 ),
    .Y(\heichips25_can_lehmann_fsm/_0208_ ),
    .B1(\heichips25_can_lehmann_fsm/_0774_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2618_  (.B1(\heichips25_can_lehmann_fsm/net485 ),
    .Y(\heichips25_can_lehmann_fsm/_0775_ ),
    .A1(\heichips25_can_lehmann_fsm/net984 ),
    .A2(\heichips25_can_lehmann_fsm/net417 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2619_  (.A1(\heichips25_can_lehmann_fsm/_0893_ ),
    .A2(\heichips25_can_lehmann_fsm/net417 ),
    .Y(\heichips25_can_lehmann_fsm/_0209_ ),
    .B1(\heichips25_can_lehmann_fsm/_0775_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2620_  (.B1(\heichips25_can_lehmann_fsm/net484 ),
    .Y(\heichips25_can_lehmann_fsm/_0776_ ),
    .A1(\heichips25_can_lehmann_fsm/net984 ),
    .A2(\heichips25_can_lehmann_fsm/net375 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2621_  (.A1(\heichips25_can_lehmann_fsm/_0892_ ),
    .A2(\heichips25_can_lehmann_fsm/net375 ),
    .Y(\heichips25_can_lehmann_fsm/_0210_ ),
    .B1(\heichips25_can_lehmann_fsm/_0776_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2622_  (.B1(\heichips25_can_lehmann_fsm/net484 ),
    .Y(\heichips25_can_lehmann_fsm/_0777_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[152] ),
    .A2(\heichips25_can_lehmann_fsm/net416 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2623_  (.A1(\heichips25_can_lehmann_fsm/_0892_ ),
    .A2(\heichips25_can_lehmann_fsm/net416 ),
    .Y(\heichips25_can_lehmann_fsm/_0211_ ),
    .B1(\heichips25_can_lehmann_fsm/_0777_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2624_  (.B1(\heichips25_can_lehmann_fsm/net482 ),
    .Y(\heichips25_can_lehmann_fsm/_0778_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[152] ),
    .A2(\heichips25_can_lehmann_fsm/net374 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2625_  (.A1(\heichips25_can_lehmann_fsm/_0891_ ),
    .A2(\heichips25_can_lehmann_fsm/net374 ),
    .Y(\heichips25_can_lehmann_fsm/_0212_ ),
    .B1(\heichips25_can_lehmann_fsm/_0778_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2626_  (.B1(\heichips25_can_lehmann_fsm/net478 ),
    .Y(\heichips25_can_lehmann_fsm/_0779_ ),
    .A1(\heichips25_can_lehmann_fsm/net963 ),
    .A2(\heichips25_can_lehmann_fsm/net409 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2627_  (.A1(\heichips25_can_lehmann_fsm/_0891_ ),
    .A2(\heichips25_can_lehmann_fsm/net409 ),
    .Y(\heichips25_can_lehmann_fsm/_0213_ ),
    .B1(\heichips25_can_lehmann_fsm/_0779_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2628_  (.B1(\heichips25_can_lehmann_fsm/net477 ),
    .Y(\heichips25_can_lehmann_fsm/_0780_ ),
    .A1(\heichips25_can_lehmann_fsm/net963 ),
    .A2(\heichips25_can_lehmann_fsm/net368 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2629_  (.A1(\heichips25_can_lehmann_fsm/_0890_ ),
    .A2(\heichips25_can_lehmann_fsm/net368 ),
    .Y(\heichips25_can_lehmann_fsm/_0214_ ),
    .B1(\heichips25_can_lehmann_fsm/_0780_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2630_  (.B1(\heichips25_can_lehmann_fsm/net476 ),
    .Y(\heichips25_can_lehmann_fsm/_0781_ ),
    .A1(\heichips25_can_lehmann_fsm/net1053 ),
    .A2(\heichips25_can_lehmann_fsm/net395 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2631_  (.A1(\heichips25_can_lehmann_fsm/_0890_ ),
    .A2(\heichips25_can_lehmann_fsm/net395 ),
    .Y(\heichips25_can_lehmann_fsm/_0215_ ),
    .B1(\heichips25_can_lehmann_fsm/_0781_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2632_  (.B1(\heichips25_can_lehmann_fsm/net479 ),
    .Y(\heichips25_can_lehmann_fsm/_0782_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[156] ),
    .A2(\heichips25_can_lehmann_fsm/net361 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2633_  (.A1(\heichips25_can_lehmann_fsm/_0889_ ),
    .A2(\heichips25_can_lehmann_fsm/net361 ),
    .Y(\heichips25_can_lehmann_fsm/_0216_ ),
    .B1(\heichips25_can_lehmann_fsm/_0782_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2634_  (.B1(\heichips25_can_lehmann_fsm/net465 ),
    .Y(\heichips25_can_lehmann_fsm/_0783_ ),
    .A1(\heichips25_can_lehmann_fsm/net964 ),
    .A2(\heichips25_can_lehmann_fsm/net394 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2635_  (.A1(\heichips25_can_lehmann_fsm/_0889_ ),
    .A2(\heichips25_can_lehmann_fsm/net394 ),
    .Y(\heichips25_can_lehmann_fsm/_0217_ ),
    .B1(\heichips25_can_lehmann_fsm/_0783_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2636_  (.B1(\heichips25_can_lehmann_fsm/net465 ),
    .Y(\heichips25_can_lehmann_fsm/_0784_ ),
    .A1(\heichips25_can_lehmann_fsm/net964 ),
    .A2(\heichips25_can_lehmann_fsm/net357 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2637_  (.A1(\heichips25_can_lehmann_fsm/_0888_ ),
    .A2(\heichips25_can_lehmann_fsm/net357 ),
    .Y(\heichips25_can_lehmann_fsm/_0218_ ),
    .B1(\heichips25_can_lehmann_fsm/_0784_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2638_  (.B1(\heichips25_can_lehmann_fsm/net468 ),
    .Y(\heichips25_can_lehmann_fsm/_0785_ ),
    .A1(\heichips25_can_lehmann_fsm/net1010 ),
    .A2(\heichips25_can_lehmann_fsm/net398 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2639_  (.A1(\heichips25_can_lehmann_fsm/_0888_ ),
    .A2(\heichips25_can_lehmann_fsm/net398 ),
    .Y(\heichips25_can_lehmann_fsm/_0219_ ),
    .B1(\heichips25_can_lehmann_fsm/_0785_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2640_  (.B1(\heichips25_can_lehmann_fsm/net468 ),
    .Y(\heichips25_can_lehmann_fsm/_0786_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[160] ),
    .A2(\heichips25_can_lehmann_fsm/net359 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2641_  (.A1(\heichips25_can_lehmann_fsm/_0887_ ),
    .A2(\heichips25_can_lehmann_fsm/net360 ),
    .Y(\heichips25_can_lehmann_fsm/_0220_ ),
    .B1(\heichips25_can_lehmann_fsm/_0786_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2642_  (.B1(\heichips25_can_lehmann_fsm/net469 ),
    .Y(\heichips25_can_lehmann_fsm/_0787_ ),
    .A1(\heichips25_can_lehmann_fsm/net1090 ),
    .A2(\heichips25_can_lehmann_fsm/net399 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2643_  (.A1(\heichips25_can_lehmann_fsm/_0887_ ),
    .A2(\heichips25_can_lehmann_fsm/net399 ),
    .Y(\heichips25_can_lehmann_fsm/_0221_ ),
    .B1(\heichips25_can_lehmann_fsm/_0787_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2644_  (.B1(\heichips25_can_lehmann_fsm/net473 ),
    .Y(\heichips25_can_lehmann_fsm/_0788_ ),
    .A1(\heichips25_can_lehmann_fsm/net855 ),
    .A2(\heichips25_can_lehmann_fsm/net401 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2645_  (.A1(\heichips25_can_lehmann_fsm/_0886_ ),
    .A2(\heichips25_can_lehmann_fsm/net401 ),
    .Y(\heichips25_can_lehmann_fsm/_0222_ ),
    .B1(\heichips25_can_lehmann_fsm/_0788_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2646_  (.B1(\heichips25_can_lehmann_fsm/net472 ),
    .Y(\heichips25_can_lehmann_fsm/_0789_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[164] ),
    .A2(\heichips25_can_lehmann_fsm/net404 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2647_  (.A1(\heichips25_can_lehmann_fsm/_0885_ ),
    .A2(\heichips25_can_lehmann_fsm/net404 ),
    .Y(\heichips25_can_lehmann_fsm/_0223_ ),
    .B1(\heichips25_can_lehmann_fsm/_0789_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2648_  (.B1(\heichips25_can_lehmann_fsm/net472 ),
    .Y(\heichips25_can_lehmann_fsm/_0790_ ),
    .A1(\heichips25_can_lehmann_fsm/net844 ),
    .A2(\heichips25_can_lehmann_fsm/net404 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2649_  (.A1(\heichips25_can_lehmann_fsm/_0884_ ),
    .A2(\heichips25_can_lehmann_fsm/net404 ),
    .Y(\heichips25_can_lehmann_fsm/_0224_ ),
    .B1(\heichips25_can_lehmann_fsm/_0790_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2650_  (.B1(\heichips25_can_lehmann_fsm/net491 ),
    .Y(\heichips25_can_lehmann_fsm/_0791_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[166] ),
    .A2(\heichips25_can_lehmann_fsm/net421 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2651_  (.A1(\heichips25_can_lehmann_fsm/_0883_ ),
    .A2(\heichips25_can_lehmann_fsm/net421 ),
    .Y(\heichips25_can_lehmann_fsm/_0225_ ),
    .B1(\heichips25_can_lehmann_fsm/_0791_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2652_  (.B1(\heichips25_can_lehmann_fsm/net492 ),
    .Y(\heichips25_can_lehmann_fsm/_0792_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[166] ),
    .A2(\heichips25_can_lehmann_fsm/net381 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2653_  (.A1(\heichips25_can_lehmann_fsm/_0882_ ),
    .A2(\heichips25_can_lehmann_fsm/net381 ),
    .Y(\heichips25_can_lehmann_fsm/_0226_ ),
    .B1(\heichips25_can_lehmann_fsm/_0792_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2654_  (.B1(\heichips25_can_lehmann_fsm/net497 ),
    .Y(\heichips25_can_lehmann_fsm/_0793_ ),
    .A1(\heichips25_can_lehmann_fsm/net1134 ),
    .A2(\heichips25_can_lehmann_fsm/net427 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2655_  (.A1(\heichips25_can_lehmann_fsm/_0882_ ),
    .A2(\heichips25_can_lehmann_fsm/net427 ),
    .Y(\heichips25_can_lehmann_fsm/_0227_ ),
    .B1(\heichips25_can_lehmann_fsm/_0793_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2656_  (.B1(\heichips25_can_lehmann_fsm/net497 ),
    .Y(\heichips25_can_lehmann_fsm/_0794_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[168] ),
    .A2(\heichips25_can_lehmann_fsm/net385 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2657_  (.A1(\heichips25_can_lehmann_fsm/_0881_ ),
    .A2(\heichips25_can_lehmann_fsm/net385 ),
    .Y(\heichips25_can_lehmann_fsm/_0228_ ),
    .B1(\heichips25_can_lehmann_fsm/_0794_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2658_  (.B1(\heichips25_can_lehmann_fsm/net497 ),
    .Y(\heichips25_can_lehmann_fsm/_0795_ ),
    .A1(\heichips25_can_lehmann_fsm/net920 ),
    .A2(\heichips25_can_lehmann_fsm/net428 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2659_  (.A1(\heichips25_can_lehmann_fsm/_0881_ ),
    .A2(\heichips25_can_lehmann_fsm/net428 ),
    .Y(\heichips25_can_lehmann_fsm/_0229_ ),
    .B1(\heichips25_can_lehmann_fsm/_0795_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2660_  (.B1(\heichips25_can_lehmann_fsm/net498 ),
    .Y(\heichips25_can_lehmann_fsm/_0796_ ),
    .A1(\heichips25_can_lehmann_fsm/net920 ),
    .A2(\heichips25_can_lehmann_fsm/net384 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2661_  (.A1(\heichips25_can_lehmann_fsm/_0880_ ),
    .A2(\heichips25_can_lehmann_fsm/net384 ),
    .Y(\heichips25_can_lehmann_fsm/_0230_ ),
    .B1(\heichips25_can_lehmann_fsm/_0796_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2662_  (.B1(\heichips25_can_lehmann_fsm/net488 ),
    .Y(\heichips25_can_lehmann_fsm/_0797_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[172] ),
    .A2(\heichips25_can_lehmann_fsm/net418 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2663_  (.A1(\heichips25_can_lehmann_fsm/_0880_ ),
    .A2(\heichips25_can_lehmann_fsm/net418 ),
    .Y(\heichips25_can_lehmann_fsm/_0231_ ),
    .B1(\heichips25_can_lehmann_fsm/_0797_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2664_  (.B1(\heichips25_can_lehmann_fsm/net487 ),
    .Y(\heichips25_can_lehmann_fsm/_0798_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[172] ),
    .A2(\heichips25_can_lehmann_fsm/net376 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2665_  (.A1(\heichips25_can_lehmann_fsm/_0879_ ),
    .A2(\heichips25_can_lehmann_fsm/net376 ),
    .Y(\heichips25_can_lehmann_fsm/_0232_ ),
    .B1(\heichips25_can_lehmann_fsm/_0798_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2666_  (.B1(\heichips25_can_lehmann_fsm/net483 ),
    .Y(\heichips25_can_lehmann_fsm/_0799_ ),
    .A1(\heichips25_can_lehmann_fsm/net1150 ),
    .A2(\heichips25_can_lehmann_fsm/net415 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2667_  (.A1(\heichips25_can_lehmann_fsm/_0879_ ),
    .A2(\heichips25_can_lehmann_fsm/net415 ),
    .Y(\heichips25_can_lehmann_fsm/_0233_ ),
    .B1(\heichips25_can_lehmann_fsm/_0799_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2668_  (.B1(\heichips25_can_lehmann_fsm/net483 ),
    .Y(\heichips25_can_lehmann_fsm/_0800_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[174] ),
    .A2(\heichips25_can_lehmann_fsm/net375 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2669_  (.A1(\heichips25_can_lehmann_fsm/_0878_ ),
    .A2(\heichips25_can_lehmann_fsm/net375 ),
    .Y(\heichips25_can_lehmann_fsm/_0234_ ),
    .B1(\heichips25_can_lehmann_fsm/_0800_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2670_  (.B1(\heichips25_can_lehmann_fsm/net484 ),
    .Y(\heichips25_can_lehmann_fsm/_0801_ ),
    .A1(\heichips25_can_lehmann_fsm/net915 ),
    .A2(\heichips25_can_lehmann_fsm/net420 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2671_  (.A1(\heichips25_can_lehmann_fsm/_0878_ ),
    .A2(\heichips25_can_lehmann_fsm/net416 ),
    .Y(\heichips25_can_lehmann_fsm/_0235_ ),
    .B1(\heichips25_can_lehmann_fsm/_0801_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2672_  (.B1(\heichips25_can_lehmann_fsm/net482 ),
    .Y(\heichips25_can_lehmann_fsm/_0802_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[176] ),
    .A2(\heichips25_can_lehmann_fsm/net374 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2673_  (.A1(\heichips25_can_lehmann_fsm/_0877_ ),
    .A2(\heichips25_can_lehmann_fsm/net374 ),
    .Y(\heichips25_can_lehmann_fsm/_0236_ ),
    .B1(\heichips25_can_lehmann_fsm/_0802_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2674_  (.B1(\heichips25_can_lehmann_fsm/net482 ),
    .Y(\heichips25_can_lehmann_fsm/_0803_ ),
    .A1(\heichips25_can_lehmann_fsm/net923 ),
    .A2(\heichips25_can_lehmann_fsm/net416 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2675_  (.A1(\heichips25_can_lehmann_fsm/_0877_ ),
    .A2(\heichips25_can_lehmann_fsm/net416 ),
    .Y(\heichips25_can_lehmann_fsm/_0237_ ),
    .B1(\heichips25_can_lehmann_fsm/_0803_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2676_  (.B1(\heichips25_can_lehmann_fsm/net477 ),
    .Y(\heichips25_can_lehmann_fsm/_0804_ ),
    .A1(\heichips25_can_lehmann_fsm/net923 ),
    .A2(\heichips25_can_lehmann_fsm/net369 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2677_  (.A1(\heichips25_can_lehmann_fsm/_0876_ ),
    .A2(\heichips25_can_lehmann_fsm/net369 ),
    .Y(\heichips25_can_lehmann_fsm/_0238_ ),
    .B1(\heichips25_can_lehmann_fsm/_0804_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2678_  (.B1(\heichips25_can_lehmann_fsm/net464 ),
    .Y(\heichips25_can_lehmann_fsm/_0805_ ),
    .A1(\heichips25_can_lehmann_fsm/net924 ),
    .A2(\heichips25_can_lehmann_fsm/net394 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2679_  (.A1(\heichips25_can_lehmann_fsm/_0876_ ),
    .A2(\heichips25_can_lehmann_fsm/net395 ),
    .Y(\heichips25_can_lehmann_fsm/_0239_ ),
    .B1(\heichips25_can_lehmann_fsm/_0805_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2680_  (.B1(\heichips25_can_lehmann_fsm/net464 ),
    .Y(\heichips25_can_lehmann_fsm/_0806_ ),
    .A1(\heichips25_can_lehmann_fsm/net924 ),
    .A2(\heichips25_can_lehmann_fsm/net357 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2681_  (.A1(\heichips25_can_lehmann_fsm/_0875_ ),
    .A2(\heichips25_can_lehmann_fsm/net358 ),
    .Y(\heichips25_can_lehmann_fsm/_0240_ ),
    .B1(\heichips25_can_lehmann_fsm/_0806_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2682_  (.B1(\heichips25_can_lehmann_fsm/net465 ),
    .Y(\heichips25_can_lehmann_fsm/_0807_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[182] ),
    .A2(\heichips25_can_lehmann_fsm/net397 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2683_  (.A1(\heichips25_can_lehmann_fsm/_0875_ ),
    .A2(\heichips25_can_lehmann_fsm/net397 ),
    .Y(\heichips25_can_lehmann_fsm/_0241_ ),
    .B1(\heichips25_can_lehmann_fsm/_0807_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2684_  (.B1(\heichips25_can_lehmann_fsm/net465 ),
    .Y(\heichips25_can_lehmann_fsm/_0808_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[182] ),
    .A2(\heichips25_can_lehmann_fsm/net358 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2685_  (.A1(\heichips25_can_lehmann_fsm/_0874_ ),
    .A2(\heichips25_can_lehmann_fsm/net359 ),
    .Y(\heichips25_can_lehmann_fsm/_0242_ ),
    .B1(\heichips25_can_lehmann_fsm/_0808_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2686_  (.B1(\heichips25_can_lehmann_fsm/net468 ),
    .Y(\heichips25_can_lehmann_fsm/_0809_ ),
    .A1(\heichips25_can_lehmann_fsm/net1033 ),
    .A2(\heichips25_can_lehmann_fsm/net398 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2687_  (.A1(\heichips25_can_lehmann_fsm/_0874_ ),
    .A2(\heichips25_can_lehmann_fsm/net398 ),
    .Y(\heichips25_can_lehmann_fsm/_0243_ ),
    .B1(\heichips25_can_lehmann_fsm/_0809_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2688_  (.B1(\heichips25_can_lehmann_fsm/net468 ),
    .Y(\heichips25_can_lehmann_fsm/_0810_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[184] ),
    .A2(\heichips25_can_lehmann_fsm/net359 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2689_  (.A1(\heichips25_can_lehmann_fsm/_0873_ ),
    .A2(\heichips25_can_lehmann_fsm/net362 ),
    .Y(\heichips25_can_lehmann_fsm/_0244_ ),
    .B1(\heichips25_can_lehmann_fsm/_0810_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2690_  (.B1(\heichips25_can_lehmann_fsm/net469 ),
    .Y(\heichips25_can_lehmann_fsm/_0811_ ),
    .A1(\heichips25_can_lehmann_fsm/net1087 ),
    .A2(\heichips25_can_lehmann_fsm/net392 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2691_  (.A1(\heichips25_can_lehmann_fsm/_0873_ ),
    .A2(\heichips25_can_lehmann_fsm/net392 ),
    .Y(\heichips25_can_lehmann_fsm/_0245_ ),
    .B1(\heichips25_can_lehmann_fsm/_0811_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2692_  (.B1(\heichips25_can_lehmann_fsm/net473 ),
    .Y(\heichips25_can_lehmann_fsm/_0812_ ),
    .A1(\heichips25_can_lehmann_fsm/net1087 ),
    .A2(\heichips25_can_lehmann_fsm/net364 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2693_  (.A1(\heichips25_can_lehmann_fsm/_0872_ ),
    .A2(\heichips25_can_lehmann_fsm/net365 ),
    .Y(\heichips25_can_lehmann_fsm/_0246_ ),
    .B1(\heichips25_can_lehmann_fsm/_0812_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2694_  (.B1(\heichips25_can_lehmann_fsm/net472 ),
    .Y(\heichips25_can_lehmann_fsm/_0813_ ),
    .A1(\heichips25_can_lehmann_fsm/net849 ),
    .A2(\heichips25_can_lehmann_fsm/net404 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2695_  (.A1(\heichips25_can_lehmann_fsm/_0872_ ),
    .A2(\heichips25_can_lehmann_fsm/net404 ),
    .Y(\heichips25_can_lehmann_fsm/_0247_ ),
    .B1(\heichips25_can_lehmann_fsm/_0813_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2696_  (.B1(\heichips25_can_lehmann_fsm/net475 ),
    .Y(\heichips25_can_lehmann_fsm/_0814_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[189] ),
    .A2(\heichips25_can_lehmann_fsm/net406 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2697_  (.A1(\heichips25_can_lehmann_fsm/_0871_ ),
    .A2(\heichips25_can_lehmann_fsm/net406 ),
    .Y(\heichips25_can_lehmann_fsm/_0248_ ),
    .B1(\heichips25_can_lehmann_fsm/_0814_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2698_  (.B1(\heichips25_can_lehmann_fsm/net494 ),
    .Y(\heichips25_can_lehmann_fsm/_0815_ ),
    .A1(\heichips25_can_lehmann_fsm/net1114 ),
    .A2(\heichips25_can_lehmann_fsm/net382 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2699_  (.A1(\heichips25_can_lehmann_fsm/_0870_ ),
    .A2(\heichips25_can_lehmann_fsm/net382 ),
    .Y(\heichips25_can_lehmann_fsm/_0249_ ),
    .B1(\heichips25_can_lehmann_fsm/_0815_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2700_  (.B1(\heichips25_can_lehmann_fsm/net495 ),
    .Y(\heichips25_can_lehmann_fsm/_0816_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[191] ),
    .A2(\heichips25_can_lehmann_fsm/net424 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2701_  (.A1(\heichips25_can_lehmann_fsm/_0870_ ),
    .A2(\heichips25_can_lehmann_fsm/net424 ),
    .Y(\heichips25_can_lehmann_fsm/_0250_ ),
    .B1(\heichips25_can_lehmann_fsm/_0816_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2702_  (.B1(\heichips25_can_lehmann_fsm/net497 ),
    .Y(\heichips25_can_lehmann_fsm/_0817_ ),
    .A1(\heichips25_can_lehmann_fsm/net1076 ),
    .A2(\heichips25_can_lehmann_fsm/net385 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2703_  (.A1(\heichips25_can_lehmann_fsm/_0869_ ),
    .A2(\heichips25_can_lehmann_fsm/net385 ),
    .Y(\heichips25_can_lehmann_fsm/_0251_ ),
    .B1(\heichips25_can_lehmann_fsm/_0817_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2704_  (.B1(\heichips25_can_lehmann_fsm/net497 ),
    .Y(\heichips25_can_lehmann_fsm/_0818_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[193] ),
    .A2(\heichips25_can_lehmann_fsm/net428 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2705_  (.A1(\heichips25_can_lehmann_fsm/_0869_ ),
    .A2(\heichips25_can_lehmann_fsm/net428 ),
    .Y(\heichips25_can_lehmann_fsm/_0252_ ),
    .B1(\heichips25_can_lehmann_fsm/_0818_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2706_  (.B1(\heichips25_can_lehmann_fsm/net502 ),
    .Y(\heichips25_can_lehmann_fsm/_0819_ ),
    .A1(\heichips25_can_lehmann_fsm/net1153 ),
    .A2(\heichips25_can_lehmann_fsm/net385 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2707_  (.A1(\heichips25_can_lehmann_fsm/_0868_ ),
    .A2(\heichips25_can_lehmann_fsm/net384 ),
    .Y(\heichips25_can_lehmann_fsm/_0253_ ),
    .B1(\heichips25_can_lehmann_fsm/_0819_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2708_  (.B1(\heichips25_can_lehmann_fsm/net486 ),
    .Y(\heichips25_can_lehmann_fsm/_0820_ ),
    .A1(\heichips25_can_lehmann_fsm/net1029 ),
    .A2(\heichips25_can_lehmann_fsm/net419 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2709_  (.A1(\heichips25_can_lehmann_fsm/_0868_ ),
    .A2(\heichips25_can_lehmann_fsm/net419 ),
    .Y(\heichips25_can_lehmann_fsm/_0254_ ),
    .B1(\heichips25_can_lehmann_fsm/_0820_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2710_  (.B1(\heichips25_can_lehmann_fsm/net486 ),
    .Y(\heichips25_can_lehmann_fsm/_0821_ ),
    .A1(\heichips25_can_lehmann_fsm/net1029 ),
    .A2(\heichips25_can_lehmann_fsm/net378 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2711_  (.A1(\heichips25_can_lehmann_fsm/_0867_ ),
    .A2(\heichips25_can_lehmann_fsm/net378 ),
    .Y(\heichips25_can_lehmann_fsm/_0255_ ),
    .B1(\heichips25_can_lehmann_fsm/_0821_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2712_  (.B1(\heichips25_can_lehmann_fsm/net485 ),
    .Y(\heichips25_can_lehmann_fsm/_0822_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[197] ),
    .A2(\heichips25_can_lehmann_fsm/net417 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2713_  (.A1(\heichips25_can_lehmann_fsm/_0867_ ),
    .A2(\heichips25_can_lehmann_fsm/net417 ),
    .Y(\heichips25_can_lehmann_fsm/_0256_ ),
    .B1(\heichips25_can_lehmann_fsm/_0822_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2714_  (.B1(\heichips25_can_lehmann_fsm/net485 ),
    .Y(\heichips25_can_lehmann_fsm/_0823_ ),
    .A1(\heichips25_can_lehmann_fsm/net1039 ),
    .A2(\heichips25_can_lehmann_fsm/net378 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2715_  (.A1(\heichips25_can_lehmann_fsm/_0866_ ),
    .A2(\heichips25_can_lehmann_fsm/net378 ),
    .Y(\heichips25_can_lehmann_fsm/_0257_ ),
    .B1(\heichips25_can_lehmann_fsm/_0823_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2716_  (.B1(\heichips25_can_lehmann_fsm/net484 ),
    .Y(\heichips25_can_lehmann_fsm/_0824_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[199] ),
    .A2(\heichips25_can_lehmann_fsm/net411 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2717_  (.A1(\heichips25_can_lehmann_fsm/_0866_ ),
    .A2(\heichips25_can_lehmann_fsm/net412 ),
    .Y(\heichips25_can_lehmann_fsm/_0258_ ),
    .B1(\heichips25_can_lehmann_fsm/_0824_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2718_  (.B1(\heichips25_can_lehmann_fsm/net478 ),
    .Y(\heichips25_can_lehmann_fsm/_0825_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[199] ),
    .A2(\heichips25_can_lehmann_fsm/net371 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2719_  (.A1(\heichips25_can_lehmann_fsm/_0865_ ),
    .A2(\heichips25_can_lehmann_fsm/net371 ),
    .Y(\heichips25_can_lehmann_fsm/_0259_ ),
    .B1(\heichips25_can_lehmann_fsm/_0825_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2720_  (.B1(\heichips25_can_lehmann_fsm/net478 ),
    .Y(\heichips25_can_lehmann_fsm/_0826_ ),
    .A1(\heichips25_can_lehmann_fsm/net1172 ),
    .A2(\heichips25_can_lehmann_fsm/net410 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2721_  (.A1(\heichips25_can_lehmann_fsm/_0865_ ),
    .A2(\heichips25_can_lehmann_fsm/net410 ),
    .Y(\heichips25_can_lehmann_fsm/_0260_ ),
    .B1(\heichips25_can_lehmann_fsm/_0826_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2722_  (.B1(\heichips25_can_lehmann_fsm/net478 ),
    .Y(\heichips25_can_lehmann_fsm/_0827_ ),
    .A1(\heichips25_can_lehmann_fsm/net1172 ),
    .A2(\heichips25_can_lehmann_fsm/net369 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2723_  (.A1(\heichips25_can_lehmann_fsm/_0864_ ),
    .A2(\heichips25_can_lehmann_fsm/net369 ),
    .Y(\heichips25_can_lehmann_fsm/_0261_ ),
    .B1(\heichips25_can_lehmann_fsm/_0827_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2724_  (.B1(\heichips25_can_lehmann_fsm/net479 ),
    .Y(\heichips25_can_lehmann_fsm/_0828_ ),
    .A1(\heichips25_can_lehmann_fsm/net848 ),
    .A2(\heichips25_can_lehmann_fsm/net410 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2725_  (.A1(\heichips25_can_lehmann_fsm/_0864_ ),
    .A2(\heichips25_can_lehmann_fsm/net410 ),
    .Y(\heichips25_can_lehmann_fsm/_0262_ ),
    .B1(\heichips25_can_lehmann_fsm/_0828_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2726_  (.B1(\heichips25_can_lehmann_fsm/net479 ),
    .Y(\heichips25_can_lehmann_fsm/_0829_ ),
    .A1(\heichips25_can_lehmann_fsm/net848 ),
    .A2(\heichips25_can_lehmann_fsm/net369 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2727_  (.A1(\heichips25_can_lehmann_fsm/_0863_ ),
    .A2(\heichips25_can_lehmann_fsm/net361 ),
    .Y(\heichips25_can_lehmann_fsm/_0263_ ),
    .B1(\heichips25_can_lehmann_fsm/_0829_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2728_  (.B1(\heichips25_can_lehmann_fsm/net465 ),
    .Y(\heichips25_can_lehmann_fsm/_0830_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[5] ),
    .A2(\heichips25_can_lehmann_fsm/net396 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2729_  (.A1(\heichips25_can_lehmann_fsm/_0863_ ),
    .A2(\heichips25_can_lehmann_fsm/net396 ),
    .Y(\heichips25_can_lehmann_fsm/_0264_ ),
    .B1(\heichips25_can_lehmann_fsm/_0830_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2730_  (.B1(\heichips25_can_lehmann_fsm/net466 ),
    .Y(\heichips25_can_lehmann_fsm/_0831_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[5] ),
    .A2(\heichips25_can_lehmann_fsm/net356 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2731_  (.A1(\heichips25_can_lehmann_fsm/_0862_ ),
    .A2(\heichips25_can_lehmann_fsm/net356 ),
    .Y(\heichips25_can_lehmann_fsm/_0265_ ),
    .B1(\heichips25_can_lehmann_fsm/_0831_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2732_  (.B1(\heichips25_can_lehmann_fsm/net466 ),
    .Y(\heichips25_can_lehmann_fsm/_0832_ ),
    .A1(\heichips25_can_lehmann_fsm/net908 ),
    .A2(\heichips25_can_lehmann_fsm/net393 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2733_  (.A1(\heichips25_can_lehmann_fsm/_0862_ ),
    .A2(\heichips25_can_lehmann_fsm/net393 ),
    .Y(\heichips25_can_lehmann_fsm/_0266_ ),
    .B1(\heichips25_can_lehmann_fsm/_0832_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2734_  (.B1(\heichips25_can_lehmann_fsm/net467 ),
    .Y(\heichips25_can_lehmann_fsm/_0833_ ),
    .A1(\heichips25_can_lehmann_fsm/net908 ),
    .A2(\heichips25_can_lehmann_fsm/net362 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2735_  (.A1(\heichips25_can_lehmann_fsm/_0861_ ),
    .A2(\heichips25_can_lehmann_fsm/net356 ),
    .Y(\heichips25_can_lehmann_fsm/_0267_ ),
    .B1(\heichips25_can_lehmann_fsm/_0833_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2736_  (.B1(\heichips25_can_lehmann_fsm/net467 ),
    .Y(\heichips25_can_lehmann_fsm/_0834_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.extended_cond.opcode[0] ),
    .A2(\heichips25_can_lehmann_fsm/net391 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2737_  (.A1(\heichips25_can_lehmann_fsm/_0861_ ),
    .A2(\heichips25_can_lehmann_fsm/net390 ),
    .Y(\heichips25_can_lehmann_fsm/_0268_ ),
    .B1(\heichips25_can_lehmann_fsm/_0834_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2738_  (.B1(\heichips25_can_lehmann_fsm/net470 ),
    .Y(\heichips25_can_lehmann_fsm/_0835_ ),
    .A1(\heichips25_can_lehmann_fsm/net343 ),
    .A2(\heichips25_can_lehmann_fsm/net355 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2739_  (.A1(\heichips25_can_lehmann_fsm/_0860_ ),
    .A2(\heichips25_can_lehmann_fsm/net355 ),
    .Y(\heichips25_can_lehmann_fsm/_0269_ ),
    .B1(\heichips25_can_lehmann_fsm/_0835_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2740_  (.B1(\heichips25_can_lehmann_fsm/net470 ),
    .Y(\heichips25_can_lehmann_fsm/_0836_ ),
    .A1(\heichips25_can_lehmann_fsm/net1154 ),
    .A2(\heichips25_can_lehmann_fsm/net391 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2741_  (.A1(\heichips25_can_lehmann_fsm/_0860_ ),
    .A2(\heichips25_can_lehmann_fsm/net391 ),
    .Y(\heichips25_can_lehmann_fsm/_0270_ ),
    .B1(\heichips25_can_lehmann_fsm/_0836_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2742_  (.B1(\heichips25_can_lehmann_fsm/net472 ),
    .Y(\heichips25_can_lehmann_fsm/_0837_ ),
    .A1(\heichips25_can_lehmann_fsm/net1154 ),
    .A2(\heichips25_can_lehmann_fsm/net365 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2743_  (.A1(\heichips25_can_lehmann_fsm/_0859_ ),
    .A2(\heichips25_can_lehmann_fsm/net365 ),
    .Y(\heichips25_can_lehmann_fsm/_0271_ ),
    .B1(\heichips25_can_lehmann_fsm/_0837_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2744_  (.B1(\heichips25_can_lehmann_fsm/net474 ),
    .Y(\heichips25_can_lehmann_fsm/_0838_ ),
    .A1(\heichips25_can_lehmann_fsm/net1147 ),
    .A2(\heichips25_can_lehmann_fsm/net405 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2745_  (.A1(\heichips25_can_lehmann_fsm/_0859_ ),
    .A2(\heichips25_can_lehmann_fsm/net405 ),
    .Y(\heichips25_can_lehmann_fsm/_0272_ ),
    .B1(\heichips25_can_lehmann_fsm/_0838_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2746_  (.B1(\heichips25_can_lehmann_fsm/net491 ),
    .Y(\heichips25_can_lehmann_fsm/_0839_ ),
    .A1(\heichips25_can_lehmann_fsm/net1127 ),
    .A2(\heichips25_can_lehmann_fsm/net421 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2747_  (.A1(\heichips25_can_lehmann_fsm/_0858_ ),
    .A2(\heichips25_can_lehmann_fsm/net421 ),
    .Y(\heichips25_can_lehmann_fsm/_0273_ ),
    .B1(\heichips25_can_lehmann_fsm/_0839_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2748_  (.B1(\heichips25_can_lehmann_fsm/net491 ),
    .Y(\heichips25_can_lehmann_fsm/_0840_ ),
    .A1(\heichips25_can_lehmann_fsm/net1127 ),
    .A2(\heichips25_can_lehmann_fsm/net380 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2749_  (.A1(\heichips25_can_lehmann_fsm/_0857_ ),
    .A2(\heichips25_can_lehmann_fsm/net381 ),
    .Y(\heichips25_can_lehmann_fsm/_0274_ ),
    .B1(\heichips25_can_lehmann_fsm/_0840_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2750_  (.B1(\heichips25_can_lehmann_fsm/net491 ),
    .Y(\heichips25_can_lehmann_fsm/_0841_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.extended_then_action[4] ),
    .A2(\heichips25_can_lehmann_fsm/net425 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2751_  (.A1(\heichips25_can_lehmann_fsm/_0857_ ),
    .A2(\heichips25_can_lehmann_fsm/net425 ),
    .Y(\heichips25_can_lehmann_fsm/_0275_ ),
    .B1(\heichips25_can_lehmann_fsm/_0841_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2752_  (.B1(\heichips25_can_lehmann_fsm/net499 ),
    .Y(\heichips25_can_lehmann_fsm/_0842_ ),
    .A1(\heichips25_can_lehmann_fsm/net1157 ),
    .A2(\heichips25_can_lehmann_fsm/net386 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2753_  (.A1(\heichips25_can_lehmann_fsm/_0856_ ),
    .A2(\heichips25_can_lehmann_fsm/net386 ),
    .Y(\heichips25_can_lehmann_fsm/_0276_ ),
    .B1(\heichips25_can_lehmann_fsm/_0842_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2754_  (.B1(\heichips25_can_lehmann_fsm/net498 ),
    .Y(\heichips25_can_lehmann_fsm/_0843_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[18] ),
    .A2(\heichips25_can_lehmann_fsm/net426 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2755_  (.A1(\heichips25_can_lehmann_fsm/_0856_ ),
    .A2(\heichips25_can_lehmann_fsm/net426 ),
    .Y(\heichips25_can_lehmann_fsm/_0277_ ),
    .B1(\heichips25_can_lehmann_fsm/_0843_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2756_  (.B1(\heichips25_can_lehmann_fsm/net498 ),
    .Y(\heichips25_can_lehmann_fsm/_0844_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[18] ),
    .A2(\heichips25_can_lehmann_fsm/net384 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2757_  (.A1(\heichips25_can_lehmann_fsm/_0855_ ),
    .A2(\heichips25_can_lehmann_fsm/net384 ),
    .Y(\heichips25_can_lehmann_fsm/_0278_ ),
    .B1(\heichips25_can_lehmann_fsm/_0844_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2758_  (.B1(\heichips25_can_lehmann_fsm/net488 ),
    .Y(\heichips25_can_lehmann_fsm/_0845_ ),
    .A1(\heichips25_can_lehmann_fsm/net1084 ),
    .A2(\heichips25_can_lehmann_fsm/net419 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2759_  (.A1(\heichips25_can_lehmann_fsm/_0855_ ),
    .A2(\heichips25_can_lehmann_fsm/net419 ),
    .Y(\heichips25_can_lehmann_fsm/_0279_ ),
    .B1(\heichips25_can_lehmann_fsm/_0845_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2760_  (.B1(\heichips25_can_lehmann_fsm/net487 ),
    .Y(\heichips25_can_lehmann_fsm/_0846_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[20] ),
    .A2(\heichips25_can_lehmann_fsm/net376 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2761_  (.A1(\heichips25_can_lehmann_fsm/_0854_ ),
    .A2(\heichips25_can_lehmann_fsm/net376 ),
    .Y(\heichips25_can_lehmann_fsm/_0280_ ),
    .B1(\heichips25_can_lehmann_fsm/_0846_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2762_  (.B1(\heichips25_can_lehmann_fsm/net487 ),
    .Y(\heichips25_can_lehmann_fsm/_0847_ ),
    .A1(\heichips25_can_lehmann_fsm/net1116 ),
    .A2(\heichips25_can_lehmann_fsm/net417 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2763_  (.A1(\heichips25_can_lehmann_fsm/_0854_ ),
    .A2(\heichips25_can_lehmann_fsm/net417 ),
    .Y(\heichips25_can_lehmann_fsm/_0281_ ),
    .B1(\heichips25_can_lehmann_fsm/_0847_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2764_  (.B1(\heichips25_can_lehmann_fsm/net487 ),
    .Y(\heichips25_can_lehmann_fsm/_0848_ ),
    .A1(\heichips25_can_lehmann_fsm/net1116 ),
    .A2(\heichips25_can_lehmann_fsm/net378 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2765_  (.A1(\heichips25_can_lehmann_fsm/_0853_ ),
    .A2(\heichips25_can_lehmann_fsm/net375 ),
    .Y(\heichips25_can_lehmann_fsm/_0282_ ),
    .B1(\heichips25_can_lehmann_fsm/_0848_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2766_  (.B1(\heichips25_can_lehmann_fsm/net485 ),
    .Y(\heichips25_can_lehmann_fsm/_0849_ ),
    .A1(\heichips25_can_lehmann_fsm/net1148 ),
    .A2(\heichips25_can_lehmann_fsm/net412 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2767_  (.A1(\heichips25_can_lehmann_fsm/_0853_ ),
    .A2(\heichips25_can_lehmann_fsm/net412 ),
    .Y(\heichips25_can_lehmann_fsm/_0283_ ),
    .B1(\heichips25_can_lehmann_fsm/_0849_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2768_  (.B1(\heichips25_can_lehmann_fsm/net480 ),
    .Y(\heichips25_can_lehmann_fsm/_0850_ ),
    .A1(\heichips25_can_lehmann_fsm/controller.extended_state[0] ),
    .A2(\heichips25_can_lehmann_fsm/net361 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2769_  (.A1(\heichips25_can_lehmann_fsm/_0852_ ),
    .A2(\heichips25_can_lehmann_fsm/net361 ),
    .Y(\heichips25_can_lehmann_fsm/_0284_ ),
    .B1(\heichips25_can_lehmann_fsm/_0850_ ));
 sg13g2_o21ai_1 \heichips25_can_lehmann_fsm/_2770_  (.B1(\heichips25_can_lehmann_fsm/net481 ),
    .Y(\heichips25_can_lehmann_fsm/_0851_ ),
    .A1(\heichips25_can_lehmann_fsm/net1137 ),
    .A2(\heichips25_can_lehmann_fsm/net400 ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2771_  (.A1(\heichips25_can_lehmann_fsm/_0852_ ),
    .A2(\heichips25_can_lehmann_fsm/net400 ),
    .Y(\heichips25_can_lehmann_fsm/_0285_ ),
    .B1(\heichips25_can_lehmann_fsm/_0851_ ));
 sg13g2_and2_1 \heichips25_can_lehmann_fsm/_2772_  (.A(\uo_out_fsm[0] ),
    .B(\heichips25_can_lehmann_fsm/net321 ),
    .X(\heichips25_can_lehmann_fsm/_0286_ ));
 sg13g2_and2_1 \heichips25_can_lehmann_fsm/_2773_  (.A(\uo_out_fsm[1] ),
    .B(\heichips25_can_lehmann_fsm/net321 ),
    .X(\heichips25_can_lehmann_fsm/_0287_ ));
 sg13g2_a21oi_1 \heichips25_can_lehmann_fsm/_2774_  (.A1(\heichips25_can_lehmann_fsm/_1041_ ),
    .A2(\heichips25_can_lehmann_fsm/_1042_ ),
    .Y(\heichips25_can_lehmann_fsm/_0288_ ),
    .B1(\heichips25_can_lehmann_fsm/_1176_ ));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2775_  (.RESET_B(net589),
    .D(\heichips25_can_lehmann_fsm/_0000_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.addr[0] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2776_  (.RESET_B(net654),
    .D(\heichips25_can_lehmann_fsm/_0001_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.addr[1] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2777_  (.RESET_B(net652),
    .D(\heichips25_can_lehmann_fsm/_0002_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.addr[2] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2778_  (.RESET_B(net650),
    .D(\heichips25_can_lehmann_fsm/net1263 ),
    .Q(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[9] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2779_  (.RESET_B(net648),
    .D(\heichips25_can_lehmann_fsm/net1254 ),
    .Q(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[10] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2780_  (.RESET_B(net646),
    .D(\heichips25_can_lehmann_fsm/net1250 ),
    .Q(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[11] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2781_  (.RESET_B(net644),
    .D(\heichips25_can_lehmann_fsm/net1261 ),
    .Q(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[12] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2782_  (.RESET_B(net642),
    .D(\heichips25_can_lehmann_fsm/net1258 ),
    .Q(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[13] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2783_  (.RESET_B(net640),
    .D(\heichips25_can_lehmann_fsm/_0008_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[14] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2784_  (.RESET_B(net638),
    .D(\heichips25_can_lehmann_fsm/net1235 ),
    .Q(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[15] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2785_  (.RESET_B(net636),
    .D(\heichips25_can_lehmann_fsm/net1252 ),
    .Q(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[16] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2786_  (.RESET_B(net634),
    .D(\heichips25_can_lehmann_fsm/net1243 ),
    .Q(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[17] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2787_  (.RESET_B(net632),
    .D(\heichips25_can_lehmann_fsm/net1241 ),
    .Q(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[18] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2788_  (.RESET_B(net630),
    .D(\heichips25_can_lehmann_fsm/_0013_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[19] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2789_  (.RESET_B(net628),
    .D(\heichips25_can_lehmann_fsm/net1247 ),
    .Q(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[20] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2790_  (.RESET_B(net626),
    .D(\heichips25_can_lehmann_fsm/net1245 ),
    .Q(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[21] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2791_  (.RESET_B(net624),
    .D(\heichips25_can_lehmann_fsm/net1239 ),
    .Q(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[22] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2792_  (.RESET_B(net622),
    .D(\heichips25_can_lehmann_fsm/net1228 ),
    .Q(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[23] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2793_  (.RESET_B(net620),
    .D(\heichips25_can_lehmann_fsm/net1256 ),
    .Q(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[8] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2794_  (.RESET_B(net618),
    .D(\heichips25_can_lehmann_fsm/_0019_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[0] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2795_  (.RESET_B(net616),
    .D(\heichips25_can_lehmann_fsm/_0020_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[1] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2796_  (.RESET_B(net614),
    .D(\heichips25_can_lehmann_fsm/_0021_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[2] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2797_  (.RESET_B(net612),
    .D(\heichips25_can_lehmann_fsm/net1220 ),
    .Q(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[3] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2798_  (.RESET_B(net610),
    .D(\heichips25_can_lehmann_fsm/net1267 ),
    .Q(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[4] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2799_  (.RESET_B(net608),
    .D(\heichips25_can_lehmann_fsm/net1265 ),
    .Q(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[5] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2800_  (.RESET_B(net606),
    .D(\heichips25_can_lehmann_fsm/net1271 ),
    .Q(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[6] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2801_  (.RESET_B(net604),
    .D(\heichips25_can_lehmann_fsm/_0026_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[7] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2802_  (.RESET_B(net602),
    .D(\heichips25_can_lehmann_fsm/_0027_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[0] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2803_  (.RESET_B(net600),
    .D(\heichips25_can_lehmann_fsm/_0028_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[1] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2804_  (.RESET_B(net598),
    .D(\heichips25_can_lehmann_fsm/net1216 ),
    .Q(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[2] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2805_  (.RESET_B(net596),
    .D(\heichips25_can_lehmann_fsm/net1203 ),
    .Q(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[3] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2806_  (.RESET_B(net594),
    .D(\heichips25_can_lehmann_fsm/net1237 ),
    .Q(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[4] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2807_  (.RESET_B(net592),
    .D(\heichips25_can_lehmann_fsm/net1211 ),
    .Q(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[5] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2808_  (.RESET_B(net590),
    .D(\heichips25_can_lehmann_fsm/net1193 ),
    .Q(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[6] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2809_  (.RESET_B(net588),
    .D(\heichips25_can_lehmann_fsm/net1199 ),
    .Q(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[7] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2810_  (.RESET_B(net586),
    .D(\heichips25_can_lehmann_fsm/_0035_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[8] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2811_  (.RESET_B(net584),
    .D(\heichips25_can_lehmann_fsm/_0036_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[9] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2812_  (.RESET_B(net582),
    .D(\heichips25_can_lehmann_fsm/net1208 ),
    .Q(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[10] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2813_  (.RESET_B(net580),
    .D(\heichips25_can_lehmann_fsm/net1187 ),
    .Q(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[11] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2814_  (.RESET_B(net578),
    .D(\heichips25_can_lehmann_fsm/net1232 ),
    .Q(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[12] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2815_  (.RESET_B(net576),
    .D(\heichips25_can_lehmann_fsm/_0040_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[13] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2816_  (.RESET_B(net574),
    .D(\heichips25_can_lehmann_fsm/net1222 ),
    .Q(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[14] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2817_  (.RESET_B(net572),
    .D(\heichips25_can_lehmann_fsm/net1206 ),
    .Q(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[15] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2818_  (.RESET_B(net570),
    .D(\heichips25_can_lehmann_fsm/_0043_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[0] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2819_  (.RESET_B(net568),
    .D(\heichips25_can_lehmann_fsm/net1175 ),
    .Q(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[1] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2820_  (.RESET_B(net566),
    .D(\heichips25_can_lehmann_fsm/net1196 ),
    .Q(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[2] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2821_  (.RESET_B(net564),
    .D(\heichips25_can_lehmann_fsm/_0046_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[3] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2822_  (.RESET_B(net562),
    .D(\heichips25_can_lehmann_fsm/net1185 ),
    .Q(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[4] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2823_  (.RESET_B(net560),
    .D(\heichips25_can_lehmann_fsm/_0048_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[5] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2824_  (.RESET_B(net558),
    .D(\heichips25_can_lehmann_fsm/_0049_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[6] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2825_  (.RESET_B(net556),
    .D(\heichips25_can_lehmann_fsm/_0050_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[7] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2826_  (.RESET_B(net554),
    .D(\heichips25_can_lehmann_fsm/_0051_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[8] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2827_  (.RESET_B(net552),
    .D(\heichips25_can_lehmann_fsm/net1171 ),
    .Q(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[9] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2828_  (.RESET_B(net550),
    .D(\heichips25_can_lehmann_fsm/_0053_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[10] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2829_  (.RESET_B(net548),
    .D(\heichips25_can_lehmann_fsm/net1166 ),
    .Q(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[11] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2830_  (.RESET_B(net546),
    .D(\heichips25_can_lehmann_fsm/_0055_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[12] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2831_  (.RESET_B(net544),
    .D(\heichips25_can_lehmann_fsm/net1159 ),
    .Q(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[13] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2832_  (.RESET_B(net542),
    .D(\heichips25_can_lehmann_fsm/net1190 ),
    .Q(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[14] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2833_  (.RESET_B(net540),
    .D(\heichips25_can_lehmann_fsm/_0058_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[15] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2834_  (.RESET_B(net538),
    .D(\heichips25_can_lehmann_fsm/_0059_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.const_data[0] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2835_  (.RESET_B(net536),
    .D(\heichips25_can_lehmann_fsm/net1094 ),
    .Q(\heichips25_can_lehmann_fsm/controller.const_data[1] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2836_  (.RESET_B(net534),
    .D(\heichips25_can_lehmann_fsm/_0061_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.const_data[2] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2837_  (.RESET_B(net532),
    .D(\heichips25_can_lehmann_fsm/net896 ),
    .Q(\heichips25_can_lehmann_fsm/controller.const_data[3] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2838_  (.RESET_B(net530),
    .D(\heichips25_can_lehmann_fsm/_0063_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.const_data[4] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2839_  (.RESET_B(net528),
    .D(\heichips25_can_lehmann_fsm/_0064_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.const_data[5] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2840_  (.RESET_B(net526),
    .D(\heichips25_can_lehmann_fsm/_0065_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.const_data[6] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2841_  (.RESET_B(net813),
    .D(\heichips25_can_lehmann_fsm/net1089 ),
    .Q(\heichips25_can_lehmann_fsm/controller.const_data[7] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2842_  (.RESET_B(net811),
    .D(\heichips25_can_lehmann_fsm/_0067_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.const_data[8] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2843_  (.RESET_B(net809),
    .D(\heichips25_can_lehmann_fsm/_0068_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.const_data[9] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2844_  (.RESET_B(net807),
    .D(\heichips25_can_lehmann_fsm/net852 ),
    .Q(\heichips25_can_lehmann_fsm/controller.const_data[10] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2845_  (.RESET_B(net805),
    .D(\heichips25_can_lehmann_fsm/net1007 ),
    .Q(\heichips25_can_lehmann_fsm/controller.const_data[11] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2846_  (.RESET_B(net803),
    .D(\heichips25_can_lehmann_fsm/_0071_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.const_data[12] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2847_  (.RESET_B(net801),
    .D(\heichips25_can_lehmann_fsm/_0072_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.const_data[13] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2848_  (.RESET_B(net799),
    .D(\heichips25_can_lehmann_fsm/_0073_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.const_data[14] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2849_  (.RESET_B(net797),
    .D(\heichips25_can_lehmann_fsm/_0074_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.const_data[15] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2850_  (.RESET_B(net795),
    .D(\heichips25_can_lehmann_fsm/_0075_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.const_data[16] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2851_  (.RESET_B(net793),
    .D(\heichips25_can_lehmann_fsm/_0076_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.const_data[17] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2852_  (.RESET_B(net791),
    .D(\heichips25_can_lehmann_fsm/net841 ),
    .Q(\heichips25_can_lehmann_fsm/controller.const_data[18] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2853_  (.RESET_B(net789),
    .D(\heichips25_can_lehmann_fsm/_0078_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.const_data[19] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2854_  (.RESET_B(net787),
    .D(\heichips25_can_lehmann_fsm/net899 ),
    .Q(\heichips25_can_lehmann_fsm/controller.const_data[20] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2855_  (.RESET_B(net785),
    .D(\heichips25_can_lehmann_fsm/net940 ),
    .Q(\heichips25_can_lehmann_fsm/controller.const_data[21] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2856_  (.RESET_B(net783),
    .D(\heichips25_can_lehmann_fsm/_0081_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.const_data[22] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2857_  (.RESET_B(net781),
    .D(\heichips25_can_lehmann_fsm/_0082_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.const_data[23] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2858_  (.RESET_B(net779),
    .D(\heichips25_can_lehmann_fsm/_0083_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.const_data[24] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2859_  (.RESET_B(net777),
    .D(\heichips25_can_lehmann_fsm/net943 ),
    .Q(\heichips25_can_lehmann_fsm/controller.const_data[25] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2860_  (.RESET_B(net775),
    .D(\heichips25_can_lehmann_fsm/_0085_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.const_data[26] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2861_  (.RESET_B(net773),
    .D(\heichips25_can_lehmann_fsm/net949 ),
    .Q(\heichips25_can_lehmann_fsm/controller.const_data[27] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2862_  (.RESET_B(net771),
    .D(\heichips25_can_lehmann_fsm/_0087_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.const_data[28] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2863_  (.RESET_B(net769),
    .D(\heichips25_can_lehmann_fsm/_0088_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.const_data[29] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2864_  (.RESET_B(net767),
    .D(\heichips25_can_lehmann_fsm/net1086 ),
    .Q(\heichips25_can_lehmann_fsm/controller.const_data[30] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2865_  (.RESET_B(net765),
    .D(\heichips25_can_lehmann_fsm/net884 ),
    .Q(\heichips25_can_lehmann_fsm/controller.const_data[31] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2866_  (.RESET_B(net763),
    .D(\heichips25_can_lehmann_fsm/_0091_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[32] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2867_  (.RESET_B(net761),
    .D(\heichips25_can_lehmann_fsm/_0092_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[33] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2868_  (.RESET_B(net759),
    .D(\heichips25_can_lehmann_fsm/_0093_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[34] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2869_  (.RESET_B(net757),
    .D(\heichips25_can_lehmann_fsm/net988 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[35] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2870_  (.RESET_B(net755),
    .D(\heichips25_can_lehmann_fsm/_0095_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[36] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2871_  (.RESET_B(net753),
    .D(\heichips25_can_lehmann_fsm/_0096_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[37] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2872_  (.RESET_B(net751),
    .D(\heichips25_can_lehmann_fsm/_0097_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[38] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2873_  (.RESET_B(net749),
    .D(\heichips25_can_lehmann_fsm/net1067 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[39] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2874_  (.RESET_B(net747),
    .D(\heichips25_can_lehmann_fsm/_0099_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[40] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2875_  (.RESET_B(net745),
    .D(\heichips25_can_lehmann_fsm/net1016 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[41] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2876_  (.RESET_B(net743),
    .D(\heichips25_can_lehmann_fsm/net1111 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[42] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2877_  (.RESET_B(net741),
    .D(\heichips25_can_lehmann_fsm/_0102_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[43] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2878_  (.RESET_B(net739),
    .D(\heichips25_can_lehmann_fsm/_0103_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[44] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2879_  (.RESET_B(net737),
    .D(\heichips25_can_lehmann_fsm/_0104_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[45] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2880_  (.RESET_B(net735),
    .D(\heichips25_can_lehmann_fsm/net1001 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[46] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2881_  (.RESET_B(net733),
    .D(\heichips25_can_lehmann_fsm/net1096 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[47] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2882_  (.RESET_B(net731),
    .D(\heichips25_can_lehmann_fsm/_0107_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[48] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2883_  (.RESET_B(net729),
    .D(\heichips25_can_lehmann_fsm/net880 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[49] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2884_  (.RESET_B(net727),
    .D(\heichips25_can_lehmann_fsm/_0109_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[50] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2885_  (.RESET_B(net725),
    .D(\heichips25_can_lehmann_fsm/_0110_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[51] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2886_  (.RESET_B(net723),
    .D(\heichips25_can_lehmann_fsm/net917 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[52] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2887_  (.RESET_B(net721),
    .D(\heichips25_can_lehmann_fsm/_0112_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[53] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2888_  (.RESET_B(net719),
    .D(\heichips25_can_lehmann_fsm/net1004 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[54] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2889_  (.RESET_B(net717),
    .D(\heichips25_can_lehmann_fsm/net871 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[55] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2890_  (.RESET_B(net715),
    .D(\heichips25_can_lehmann_fsm/_0115_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[56] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2891_  (.RESET_B(net713),
    .D(\heichips25_can_lehmann_fsm/net956 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[57] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2892_  (.RESET_B(net711),
    .D(\heichips25_can_lehmann_fsm/_0117_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[58] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2893_  (.RESET_B(net709),
    .D(\heichips25_can_lehmann_fsm/_0118_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[59] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2894_  (.RESET_B(net707),
    .D(\heichips25_can_lehmann_fsm/net1101 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[60] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2895_  (.RESET_B(net705),
    .D(\heichips25_can_lehmann_fsm/net866 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[61] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2896_  (.RESET_B(net703),
    .D(\heichips25_can_lehmann_fsm/_0121_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[62] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2897_  (.RESET_B(net701),
    .D(\heichips25_can_lehmann_fsm/_0122_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[63] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2898_  (.RESET_B(net699),
    .D(\heichips25_can_lehmann_fsm/net914 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[64] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2899_  (.RESET_B(net697),
    .D(\heichips25_can_lehmann_fsm/net1057 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[65] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2900_  (.RESET_B(net695),
    .D(\heichips25_can_lehmann_fsm/_0125_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[66] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2901_  (.RESET_B(net693),
    .D(\heichips25_can_lehmann_fsm/net1009 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[67] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2902_  (.RESET_B(net691),
    .D(\heichips25_can_lehmann_fsm/_0127_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[68] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2903_  (.RESET_B(net689),
    .D(\heichips25_can_lehmann_fsm/_0128_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[69] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2904_  (.RESET_B(net687),
    .D(\heichips25_can_lehmann_fsm/net997 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[70] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2905_  (.RESET_B(net685),
    .D(\heichips25_can_lehmann_fsm/net1042 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[71] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2906_  (.RESET_B(net683),
    .D(\heichips25_can_lehmann_fsm/_0131_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[72] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2907_  (.RESET_B(net681),
    .D(\heichips25_can_lehmann_fsm/net901 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[73] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2908_  (.RESET_B(net679),
    .D(\heichips25_can_lehmann_fsm/_0133_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[74] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2909_  (.RESET_B(net677),
    .D(\heichips25_can_lehmann_fsm/_0134_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[75] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2910_  (.RESET_B(net675),
    .D(\heichips25_can_lehmann_fsm/net910 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[76] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2911_  (.RESET_B(net673),
    .D(\heichips25_can_lehmann_fsm/net967 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[77] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2912_  (.RESET_B(net671),
    .D(\heichips25_can_lehmann_fsm/_0137_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[78] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2913_  (.RESET_B(net669),
    .D(\heichips25_can_lehmann_fsm/_0138_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[79] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2914_  (.RESET_B(net667),
    .D(\heichips25_can_lehmann_fsm/_0139_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[80] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2915_  (.RESET_B(net665),
    .D(\heichips25_can_lehmann_fsm/_0140_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[81] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2916_  (.RESET_B(net663),
    .D(\heichips25_can_lehmann_fsm/net862 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[82] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2917_  (.RESET_B(net661),
    .D(\heichips25_can_lehmann_fsm/_0142_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[83] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2918_  (.RESET_B(net659),
    .D(\heichips25_can_lehmann_fsm/_0143_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[84] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2919_  (.RESET_B(net657),
    .D(\heichips25_can_lehmann_fsm/_0144_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[85] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2920_  (.RESET_B(net655),
    .D(\heichips25_can_lehmann_fsm/net982 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[86] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2921_  (.RESET_B(net651),
    .D(\heichips25_can_lehmann_fsm/net938 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[87] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2922_  (.RESET_B(net647),
    .D(\heichips25_can_lehmann_fsm/_0147_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[88] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2923_  (.RESET_B(net643),
    .D(\heichips25_can_lehmann_fsm/_0148_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[89] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2924_  (.RESET_B(net639),
    .D(\heichips25_can_lehmann_fsm/net894 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[90] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2925_  (.RESET_B(net635),
    .D(\heichips25_can_lehmann_fsm/_0150_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[91] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2926_  (.RESET_B(net631),
    .D(\heichips25_can_lehmann_fsm/net1048 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[92] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2927_  (.RESET_B(net627),
    .D(\heichips25_can_lehmann_fsm/_0152_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[93] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2928_  (.RESET_B(net623),
    .D(\heichips25_can_lehmann_fsm/net1063 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[94] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2929_  (.RESET_B(net619),
    .D(\heichips25_can_lehmann_fsm/net859 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[95] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2930_  (.RESET_B(net615),
    .D(\heichips25_can_lehmann_fsm/_0155_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[96] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2931_  (.RESET_B(net611),
    .D(\heichips25_can_lehmann_fsm/_0156_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[97] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2932_  (.RESET_B(net607),
    .D(\heichips25_can_lehmann_fsm/_0157_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[98] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2933_  (.RESET_B(net603),
    .D(\heichips25_can_lehmann_fsm/_0158_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[99] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2934_  (.RESET_B(net599),
    .D(\heichips25_can_lehmann_fsm/net864 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[100] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2935_  (.RESET_B(net595),
    .D(\heichips25_can_lehmann_fsm/net1107 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[101] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2936_  (.RESET_B(net591),
    .D(\heichips25_can_lehmann_fsm/_0161_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[102] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2937_  (.RESET_B(net587),
    .D(\heichips25_can_lehmann_fsm/_0162_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[103] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2938_  (.RESET_B(net583),
    .D(\heichips25_can_lehmann_fsm/net1014 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[104] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2939_  (.RESET_B(net579),
    .D(\heichips25_can_lehmann_fsm/net1098 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[105] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2940_  (.RESET_B(net575),
    .D(\heichips25_can_lehmann_fsm/_0165_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[106] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2941_  (.RESET_B(net571),
    .D(\heichips25_can_lehmann_fsm/_0166_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[107] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2942_  (.RESET_B(net567),
    .D(\heichips25_can_lehmann_fsm/net971 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[108] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2943_  (.RESET_B(net563),
    .D(\heichips25_can_lehmann_fsm/net1026 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[109] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2944_  (.RESET_B(net559),
    .D(\heichips25_can_lehmann_fsm/_0169_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[110] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2945_  (.RESET_B(net555),
    .D(\heichips25_can_lehmann_fsm/_0170_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[111] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2946_  (.RESET_B(net551),
    .D(\heichips25_can_lehmann_fsm/net905 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[112] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2947_  (.RESET_B(net547),
    .D(\heichips25_can_lehmann_fsm/net935 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[113] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2948_  (.RESET_B(net543),
    .D(\heichips25_can_lehmann_fsm/_0173_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[114] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2949_  (.RESET_B(net539),
    .D(\heichips25_can_lehmann_fsm/_0174_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[115] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2950_  (.RESET_B(net535),
    .D(\heichips25_can_lehmann_fsm/net1061 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[116] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2951_  (.RESET_B(net531),
    .D(\heichips25_can_lehmann_fsm/net1078 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[117] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2952_  (.RESET_B(net527),
    .D(\heichips25_can_lehmann_fsm/_0177_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[118] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2953_  (.RESET_B(net812),
    .D(\heichips25_can_lehmann_fsm/_0178_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[119] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2954_  (.RESET_B(net808),
    .D(\heichips25_can_lehmann_fsm/net1104 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[120] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2955_  (.RESET_B(net804),
    .D(\heichips25_can_lehmann_fsm/net1028 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[121] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2956_  (.RESET_B(net800),
    .D(\heichips25_can_lehmann_fsm/_0181_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[122] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2957_  (.RESET_B(net796),
    .D(\heichips25_can_lehmann_fsm/net1036 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[123] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2958_  (.RESET_B(net792),
    .D(\heichips25_can_lehmann_fsm/_0183_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[124] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2959_  (.RESET_B(net788),
    .D(\heichips25_can_lehmann_fsm/_0184_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[125] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2960_  (.RESET_B(net784),
    .D(\heichips25_can_lehmann_fsm/net1046 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[126] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2961_  (.RESET_B(net780),
    .D(\heichips25_can_lehmann_fsm/net1018 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[127] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2962_  (.RESET_B(net776),
    .D(\heichips25_can_lehmann_fsm/_0187_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[128] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2963_  (.RESET_B(net772),
    .D(\heichips25_can_lehmann_fsm/_0188_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[129] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2964_  (.RESET_B(net768),
    .D(\heichips25_can_lehmann_fsm/_0189_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[130] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2965_  (.RESET_B(net764),
    .D(\heichips25_can_lehmann_fsm/net875 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[131] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2966_  (.RESET_B(net760),
    .D(\heichips25_can_lehmann_fsm/_0191_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[132] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2967_  (.RESET_B(net756),
    .D(\heichips25_can_lehmann_fsm/net886 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[133] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2968_  (.RESET_B(net752),
    .D(\heichips25_can_lehmann_fsm/_0193_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[134] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2969_  (.RESET_B(net748),
    .D(\heichips25_can_lehmann_fsm/_0194_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[135] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2970_  (.RESET_B(net744),
    .D(\heichips25_can_lehmann_fsm/net888 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[136] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2971_  (.RESET_B(net740),
    .D(\heichips25_can_lehmann_fsm/net947 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[137] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2972_  (.RESET_B(net736),
    .D(\heichips25_can_lehmann_fsm/_0197_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[138] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2973_  (.RESET_B(net732),
    .D(\heichips25_can_lehmann_fsm/_0198_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[139] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2974_  (.RESET_B(net728),
    .D(\heichips25_can_lehmann_fsm/net958 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[140] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2975_  (.RESET_B(net724),
    .D(\heichips25_can_lehmann_fsm/_0200_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[141] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2976_  (.RESET_B(net720),
    .D(\heichips25_can_lehmann_fsm/net847 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[142] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2977_  (.RESET_B(net716),
    .D(\heichips25_can_lehmann_fsm/_0202_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[143] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2978_  (.RESET_B(net712),
    .D(\heichips25_can_lehmann_fsm/_0203_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[144] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2979_  (.RESET_B(net708),
    .D(\heichips25_can_lehmann_fsm/_0204_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[145] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2980_  (.RESET_B(net704),
    .D(\heichips25_can_lehmann_fsm/net873 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[146] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2981_  (.RESET_B(net700),
    .D(\heichips25_can_lehmann_fsm/net1023 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[147] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2982_  (.RESET_B(net696),
    .D(\heichips25_can_lehmann_fsm/_0207_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[148] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2983_  (.RESET_B(net692),
    .D(\heichips25_can_lehmann_fsm/net986 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[149] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2984_  (.RESET_B(net688),
    .D(\heichips25_can_lehmann_fsm/_0209_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[150] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2985_  (.RESET_B(net684),
    .D(\heichips25_can_lehmann_fsm/_0210_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[151] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2986_  (.RESET_B(net680),
    .D(\heichips25_can_lehmann_fsm/net979 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[152] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2987_  (.RESET_B(net676),
    .D(\heichips25_can_lehmann_fsm/net890 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[153] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2988_  (.RESET_B(net672),
    .D(\heichips25_can_lehmann_fsm/_0213_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[154] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2989_  (.RESET_B(net668),
    .D(\heichips25_can_lehmann_fsm/_0214_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[155] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2990_  (.RESET_B(net664),
    .D(\heichips25_can_lehmann_fsm/_0215_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[156] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2991_  (.RESET_B(net660),
    .D(\heichips25_can_lehmann_fsm/net919 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[157] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2992_  (.RESET_B(net656),
    .D(\heichips25_can_lehmann_fsm/_0217_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[158] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2993_  (.RESET_B(net649),
    .D(\heichips25_can_lehmann_fsm/_0218_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[159] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2994_  (.RESET_B(net641),
    .D(\heichips25_can_lehmann_fsm/_0219_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[160] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2995_  (.RESET_B(net633),
    .D(\heichips25_can_lehmann_fsm/net929 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[161] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2996_  (.RESET_B(net625),
    .D(\heichips25_can_lehmann_fsm/_0221_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[162] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2997_  (.RESET_B(net617),
    .D(\heichips25_can_lehmann_fsm/_0222_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[163] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2998_  (.RESET_B(net609),
    .D(\heichips25_can_lehmann_fsm/net856 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[164] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_2999_  (.RESET_B(net601),
    .D(\heichips25_can_lehmann_fsm/_0224_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[165] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3000_  (.RESET_B(net593),
    .D(\heichips25_can_lehmann_fsm/net845 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[166] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3001_  (.RESET_B(net585),
    .D(\heichips25_can_lehmann_fsm/net1123 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[167] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3002_  (.RESET_B(net577),
    .D(\heichips25_can_lehmann_fsm/_0227_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[168] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3003_  (.RESET_B(net569),
    .D(\heichips25_can_lehmann_fsm/net907 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[169] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3004_  (.RESET_B(net561),
    .D(\heichips25_can_lehmann_fsm/_0229_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[170] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3005_  (.RESET_B(net553),
    .D(\heichips25_can_lehmann_fsm/_0230_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[171] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3006_  (.RESET_B(net545),
    .D(\heichips25_can_lehmann_fsm/net932 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[172] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3007_  (.RESET_B(net537),
    .D(\heichips25_can_lehmann_fsm/net1140 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[173] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3008_  (.RESET_B(net529),
    .D(\heichips25_can_lehmann_fsm/_0233_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[174] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3009_  (.RESET_B(net810),
    .D(\heichips25_can_lehmann_fsm/net868 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[175] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3010_  (.RESET_B(net802),
    .D(\heichips25_can_lehmann_fsm/_0235_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[176] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3011_  (.RESET_B(net794),
    .D(\heichips25_can_lehmann_fsm/net882 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[177] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3012_  (.RESET_B(net786),
    .D(\heichips25_can_lehmann_fsm/_0237_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[178] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3013_  (.RESET_B(net778),
    .D(\heichips25_can_lehmann_fsm/_0238_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[179] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3014_  (.RESET_B(net770),
    .D(\heichips25_can_lehmann_fsm/_0239_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[180] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3015_  (.RESET_B(net762),
    .D(\heichips25_can_lehmann_fsm/_0240_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[181] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3016_  (.RESET_B(net754),
    .D(\heichips25_can_lehmann_fsm/net854 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[182] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3017_  (.RESET_B(net746),
    .D(\heichips25_can_lehmann_fsm/net999 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[183] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3018_  (.RESET_B(net738),
    .D(\heichips25_can_lehmann_fsm/_0243_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[184] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3019_  (.RESET_B(net730),
    .D(\heichips25_can_lehmann_fsm/net991 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[185] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3020_  (.RESET_B(net722),
    .D(\heichips25_can_lehmann_fsm/_0245_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[186] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3021_  (.RESET_B(net714),
    .D(\heichips25_can_lehmann_fsm/_0246_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[187] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3022_  (.RESET_B(net706),
    .D(\heichips25_can_lehmann_fsm/_0247_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[188] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3023_  (.RESET_B(net698),
    .D(\heichips25_can_lehmann_fsm/net850 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[189] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3024_  (.RESET_B(net690),
    .D(\heichips25_can_lehmann_fsm/_0249_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[190] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3025_  (.RESET_B(net682),
    .D(\heichips25_can_lehmann_fsm/net1075 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[191] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3026_  (.RESET_B(net674),
    .D(\heichips25_can_lehmann_fsm/_0251_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[192] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3027_  (.RESET_B(net666),
    .D(\heichips25_can_lehmann_fsm/net961 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[193] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3028_  (.RESET_B(net658),
    .D(\heichips25_can_lehmann_fsm/_0253_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[194] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3029_  (.RESET_B(net645),
    .D(\heichips25_can_lehmann_fsm/_0254_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[195] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3030_  (.RESET_B(net629),
    .D(\heichips25_can_lehmann_fsm/_0255_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[196] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3031_  (.RESET_B(net613),
    .D(\heichips25_can_lehmann_fsm/net952 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[197] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3032_  (.RESET_B(net597),
    .D(\heichips25_can_lehmann_fsm/_0257_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[198] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3033_  (.RESET_B(net581),
    .D(\heichips25_can_lehmann_fsm/net994 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[199] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3034_  (.RESET_B(net565),
    .D(\heichips25_can_lehmann_fsm/net1161 ),
    .Q(\heichips25_can_lehmann_fsm/controller.extended_jump_target[0] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3035_  (.RESET_B(net549),
    .D(\heichips25_can_lehmann_fsm/_0260_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.extended_jump_target[1] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3036_  (.RESET_B(net533),
    .D(\heichips25_can_lehmann_fsm/_0261_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.extended_jump_target[2] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3037_  (.RESET_B(net806),
    .D(\heichips25_can_lehmann_fsm/_0262_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[3] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3038_  (.RESET_B(net790),
    .D(\heichips25_can_lehmann_fsm/_0263_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[4] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3039_  (.RESET_B(net774),
    .D(\heichips25_can_lehmann_fsm/net843 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[5] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3040_  (.RESET_B(net758),
    .D(\heichips25_can_lehmann_fsm/net945 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[6] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3041_  (.RESET_B(net742),
    .D(\heichips25_can_lehmann_fsm/_0266_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[7] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3042_  (.RESET_B(net726),
    .D(\heichips25_can_lehmann_fsm/_0267_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[8] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3043_  (.RESET_B(net710),
    .D(\heichips25_can_lehmann_fsm/net878 ),
    .Q(\heichips25_can_lehmann_fsm/controller.extended_cond.opcode[0] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3044_  (.RESET_B(net694),
    .D(\heichips25_can_lehmann_fsm/net1230 ),
    .Q(\heichips25_can_lehmann_fsm/controller.extended_cond.opcode[1] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3045_  (.RESET_B(net678),
    .D(\heichips25_can_lehmann_fsm/_0270_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.extended_cond.opcode[2] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3046_  (.RESET_B(net662),
    .D(\heichips25_can_lehmann_fsm/_0271_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.extended_then_action[0] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3047_  (.RESET_B(net637),
    .D(\heichips25_can_lehmann_fsm/_0272_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.extended_then_action[1] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3048_  (.RESET_B(net605),
    .D(\heichips25_can_lehmann_fsm/_0273_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.extended_then_action[2] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3049_  (.RESET_B(net573),
    .D(\heichips25_can_lehmann_fsm/_0274_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.extended_then_action[3] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3050_  (.RESET_B(net541),
    .D(\heichips25_can_lehmann_fsm/net1118 ),
    .Q(\heichips25_can_lehmann_fsm/controller.extended_then_action[4] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3051_  (.RESET_B(net798),
    .D(\heichips25_can_lehmann_fsm/_0276_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.extended_then_action[5] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3052_  (.RESET_B(net766),
    .D(\heichips25_can_lehmann_fsm/net1156 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[18] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3053_  (.RESET_B(net734),
    .D(\heichips25_can_lehmann_fsm/net1052 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[19] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3054_  (.RESET_B(net702),
    .D(\heichips25_can_lehmann_fsm/_0279_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[20] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3055_  (.RESET_B(net670),
    .D(\heichips25_can_lehmann_fsm/net1044 ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[21] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3056_  (.RESET_B(net621),
    .D(\heichips25_can_lehmann_fsm/_0281_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[22] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3057_  (.RESET_B(net557),
    .D(\heichips25_can_lehmann_fsm/_0282_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[23] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3058_  (.RESET_B(net782),
    .D(\heichips25_can_lehmann_fsm/_0283_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.extended_state[0] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3059_  (.RESET_B(net718),
    .D(\heichips25_can_lehmann_fsm/net1133 ),
    .Q(\heichips25_can_lehmann_fsm/controller.extended_state[1] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3060_  (.RESET_B(net653),
    .D(\heichips25_can_lehmann_fsm/_0285_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.extended_state[2] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3061_  (.RESET_B(net525),
    .D(\heichips25_can_lehmann_fsm/_0286_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.output_controller.keep[0] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3062_  (.RESET_B(net750),
    .D(\heichips25_can_lehmann_fsm/_0287_ ),
    .Q(\heichips25_can_lehmann_fsm/controller.output_controller.keep[1] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 \heichips25_can_lehmann_fsm/_3063_  (.RESET_B(net686),
    .D(\heichips25_can_lehmann_fsm/net1214 ),
    .Q(\heichips25_can_lehmann_fsm/controller.output_controller.keep[2] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2840__527  (.L_HI(net526));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2952__528  (.L_HI(net527));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2839__529  (.L_HI(net528));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3008__530  (.L_HI(net529));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2838__531  (.L_HI(net530));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2951__532  (.L_HI(net531));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2837__533  (.L_HI(net532));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3036__534  (.L_HI(net533));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2836__535  (.L_HI(net534));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2950__536  (.L_HI(net535));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2835__537  (.L_HI(net536));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3007__538  (.L_HI(net537));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2834__539  (.L_HI(net538));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2949__540  (.L_HI(net539));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2833__541  (.L_HI(net540));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3050__542  (.L_HI(net541));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2832__543  (.L_HI(net542));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2948__544  (.L_HI(net543));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2831__545  (.L_HI(net544));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3006__546  (.L_HI(net545));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2830__547  (.L_HI(net546));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2947__548  (.L_HI(net547));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2829__549  (.L_HI(net548));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3035__550  (.L_HI(net549));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2828__551  (.L_HI(net550));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2946__552  (.L_HI(net551));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2827__553  (.L_HI(net552));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3005__554  (.L_HI(net553));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2826__555  (.L_HI(net554));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2945__556  (.L_HI(net555));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2825__557  (.L_HI(net556));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3057__558  (.L_HI(net557));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2824__559  (.L_HI(net558));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2944__560  (.L_HI(net559));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2823__561  (.L_HI(net560));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3004__562  (.L_HI(net561));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2822__563  (.L_HI(net562));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2943__564  (.L_HI(net563));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2821__565  (.L_HI(net564));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3034__566  (.L_HI(net565));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2820__567  (.L_HI(net566));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2942__568  (.L_HI(net567));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2819__569  (.L_HI(net568));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3003__570  (.L_HI(net569));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2818__571  (.L_HI(net570));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2941__572  (.L_HI(net571));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2817__573  (.L_HI(net572));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3049__574  (.L_HI(net573));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2816__575  (.L_HI(net574));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2940__576  (.L_HI(net575));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2815__577  (.L_HI(net576));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3002__578  (.L_HI(net577));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2814__579  (.L_HI(net578));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2939__580  (.L_HI(net579));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2813__581  (.L_HI(net580));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3033__582  (.L_HI(net581));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2812__583  (.L_HI(net582));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2938__584  (.L_HI(net583));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2811__585  (.L_HI(net584));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3001__586  (.L_HI(net585));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2810__587  (.L_HI(net586));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2937__588  (.L_HI(net587));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2809__589  (.L_HI(net588));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2775__590  (.L_HI(net589));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2808__591  (.L_HI(net590));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2936__592  (.L_HI(net591));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2807__593  (.L_HI(net592));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3000__594  (.L_HI(net593));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2806__595  (.L_HI(net594));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2935__596  (.L_HI(net595));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2805__597  (.L_HI(net596));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3032__598  (.L_HI(net597));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2804__599  (.L_HI(net598));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2934__600  (.L_HI(net599));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2803__601  (.L_HI(net600));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2999__602  (.L_HI(net601));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2802__603  (.L_HI(net602));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2933__604  (.L_HI(net603));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2801__605  (.L_HI(net604));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3048__606  (.L_HI(net605));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2800__607  (.L_HI(net606));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2932__608  (.L_HI(net607));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2799__609  (.L_HI(net608));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2998__610  (.L_HI(net609));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2798__611  (.L_HI(net610));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2931__612  (.L_HI(net611));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2797__613  (.L_HI(net612));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3031__614  (.L_HI(net613));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2796__615  (.L_HI(net614));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2930__616  (.L_HI(net615));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2795__617  (.L_HI(net616));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2997__618  (.L_HI(net617));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2794__619  (.L_HI(net618));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2929__620  (.L_HI(net619));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2793__621  (.L_HI(net620));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3056__622  (.L_HI(net621));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2792__623  (.L_HI(net622));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2928__624  (.L_HI(net623));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2791__625  (.L_HI(net624));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2996__626  (.L_HI(net625));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2790__627  (.L_HI(net626));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2927__628  (.L_HI(net627));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2789__629  (.L_HI(net628));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3030__630  (.L_HI(net629));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2788__631  (.L_HI(net630));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2926__632  (.L_HI(net631));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2787__633  (.L_HI(net632));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2995__634  (.L_HI(net633));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2786__635  (.L_HI(net634));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2925__636  (.L_HI(net635));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2785__637  (.L_HI(net636));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3047__638  (.L_HI(net637));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2784__639  (.L_HI(net638));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2924__640  (.L_HI(net639));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2783__641  (.L_HI(net640));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2994__642  (.L_HI(net641));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2782__643  (.L_HI(net642));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2923__644  (.L_HI(net643));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2781__645  (.L_HI(net644));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3029__646  (.L_HI(net645));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2780__647  (.L_HI(net646));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2922__648  (.L_HI(net647));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2779__649  (.L_HI(net648));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2993__650  (.L_HI(net649));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2778__651  (.L_HI(net650));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2921__652  (.L_HI(net651));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2777__653  (.L_HI(net652));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3060__654  (.L_HI(net653));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2776__655  (.L_HI(net654));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2920__656  (.L_HI(net655));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2992__657  (.L_HI(net656));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2919__658  (.L_HI(net657));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3028__659  (.L_HI(net658));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2918__660  (.L_HI(net659));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2991__661  (.L_HI(net660));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2917__662  (.L_HI(net661));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3046__663  (.L_HI(net662));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2916__664  (.L_HI(net663));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2990__665  (.L_HI(net664));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2915__666  (.L_HI(net665));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3027__667  (.L_HI(net666));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2914__668  (.L_HI(net667));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2989__669  (.L_HI(net668));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2913__670  (.L_HI(net669));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3055__671  (.L_HI(net670));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2912__672  (.L_HI(net671));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2988__673  (.L_HI(net672));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2911__674  (.L_HI(net673));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3026__675  (.L_HI(net674));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2910__676  (.L_HI(net675));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2987__677  (.L_HI(net676));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2909__678  (.L_HI(net677));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3045__679  (.L_HI(net678));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2908__680  (.L_HI(net679));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2986__681  (.L_HI(net680));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2907__682  (.L_HI(net681));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3025__683  (.L_HI(net682));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2906__684  (.L_HI(net683));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2985__685  (.L_HI(net684));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2905__686  (.L_HI(net685));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3063__687  (.L_HI(net686));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2904__688  (.L_HI(net687));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2984__689  (.L_HI(net688));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2903__690  (.L_HI(net689));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3024__691  (.L_HI(net690));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2902__692  (.L_HI(net691));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2983__693  (.L_HI(net692));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2901__694  (.L_HI(net693));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3044__695  (.L_HI(net694));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2900__696  (.L_HI(net695));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2982__697  (.L_HI(net696));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2899__698  (.L_HI(net697));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3023__699  (.L_HI(net698));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2898__700  (.L_HI(net699));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2981__701  (.L_HI(net700));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2897__702  (.L_HI(net701));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3054__703  (.L_HI(net702));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2896__704  (.L_HI(net703));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2980__705  (.L_HI(net704));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2895__706  (.L_HI(net705));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3022__707  (.L_HI(net706));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2894__708  (.L_HI(net707));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2979__709  (.L_HI(net708));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2893__710  (.L_HI(net709));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3043__711  (.L_HI(net710));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2892__712  (.L_HI(net711));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2978__713  (.L_HI(net712));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2891__714  (.L_HI(net713));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3021__715  (.L_HI(net714));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2890__716  (.L_HI(net715));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2977__717  (.L_HI(net716));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2889__718  (.L_HI(net717));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3059__719  (.L_HI(net718));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2888__720  (.L_HI(net719));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2976__721  (.L_HI(net720));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2887__722  (.L_HI(net721));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3020__723  (.L_HI(net722));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2886__724  (.L_HI(net723));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2975__725  (.L_HI(net724));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2885__726  (.L_HI(net725));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3042__727  (.L_HI(net726));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2884__728  (.L_HI(net727));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2974__729  (.L_HI(net728));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2883__730  (.L_HI(net729));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3019__731  (.L_HI(net730));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2882__732  (.L_HI(net731));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2973__733  (.L_HI(net732));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2881__734  (.L_HI(net733));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3053__735  (.L_HI(net734));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2880__736  (.L_HI(net735));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2972__737  (.L_HI(net736));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2879__738  (.L_HI(net737));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3018__739  (.L_HI(net738));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2878__740  (.L_HI(net739));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2971__741  (.L_HI(net740));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2877__742  (.L_HI(net741));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3041__743  (.L_HI(net742));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2876__744  (.L_HI(net743));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2970__745  (.L_HI(net744));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2875__746  (.L_HI(net745));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3017__747  (.L_HI(net746));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2874__748  (.L_HI(net747));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2969__749  (.L_HI(net748));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2873__750  (.L_HI(net749));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3062__751  (.L_HI(net750));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2872__752  (.L_HI(net751));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2968__753  (.L_HI(net752));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2871__754  (.L_HI(net753));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3016__755  (.L_HI(net754));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2870__756  (.L_HI(net755));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2967__757  (.L_HI(net756));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2869__758  (.L_HI(net757));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3040__759  (.L_HI(net758));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2868__760  (.L_HI(net759));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2966__761  (.L_HI(net760));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2867__762  (.L_HI(net761));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3015__763  (.L_HI(net762));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2866__764  (.L_HI(net763));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2965__765  (.L_HI(net764));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2865__766  (.L_HI(net765));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3052__767  (.L_HI(net766));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2864__768  (.L_HI(net767));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2964__769  (.L_HI(net768));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2863__770  (.L_HI(net769));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3014__771  (.L_HI(net770));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2862__772  (.L_HI(net771));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2963__773  (.L_HI(net772));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2861__774  (.L_HI(net773));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3039__775  (.L_HI(net774));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2860__776  (.L_HI(net775));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2962__777  (.L_HI(net776));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2859__778  (.L_HI(net777));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3013__779  (.L_HI(net778));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2858__780  (.L_HI(net779));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2961__781  (.L_HI(net780));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2857__782  (.L_HI(net781));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3058__783  (.L_HI(net782));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2856__784  (.L_HI(net783));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2960__785  (.L_HI(net784));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2855__786  (.L_HI(net785));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3012__787  (.L_HI(net786));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2854__788  (.L_HI(net787));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2959__789  (.L_HI(net788));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2853__790  (.L_HI(net789));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3038__791  (.L_HI(net790));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2852__792  (.L_HI(net791));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2958__793  (.L_HI(net792));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2851__794  (.L_HI(net793));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3011__795  (.L_HI(net794));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2850__796  (.L_HI(net795));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2957__797  (.L_HI(net796));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2849__798  (.L_HI(net797));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3051__799  (.L_HI(net798));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2848__800  (.L_HI(net799));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2956__801  (.L_HI(net800));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2847__802  (.L_HI(net801));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3010__803  (.L_HI(net802));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2846__804  (.L_HI(net803));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2955__805  (.L_HI(net804));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2845__806  (.L_HI(net805));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3037__807  (.L_HI(net806));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2844__808  (.L_HI(net807));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2954__809  (.L_HI(net808));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2843__810  (.L_HI(net809));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_3009__811  (.L_HI(net810));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2842__812  (.L_HI(net811));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2953__813  (.L_HI(net812));
 sg13g2_tiehi \heichips25_can_lehmann_fsm/_2841__814  (.L_HI(net813));
 sg13g2_inv_1 \heichips25_sap3/_2003__815  (.Y(net814),
    .A(\clknet_5_24__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_tielo _23__509 (.L_LO(net508));
 sg13g2_tielo _24__510 (.L_LO(net509));
 sg13g2_tielo _25__511 (.L_LO(net510));
 sg13g2_tielo _26__512 (.L_LO(net511));
 sg13g2_tielo _27__513 (.L_LO(net512));
 sg13g2_tielo _28__514 (.L_LO(net513));
 sg13g2_tielo _29__515 (.L_LO(net514));
 sg13g2_tielo _14__516 (.L_LO(net515));
 sg13g2_tielo _15__517 (.L_LO(net516));
 sg13g2_tielo _16__518 (.L_LO(net517));
 sg13g2_tielo _17__519 (.L_LO(net518));
 sg13g2_tielo _18__520 (.L_LO(net519));
 sg13g2_tielo _19__521 (.L_LO(net520));
 sg13g2_tielo _20__522 (.L_LO(net521));
 sg13g2_tielo _21__523 (.L_LO(net522));
 sg13g2_tielo _12__524 (.L_LO(net523));
 sg13g2_inv_1 \heichips25_sap3/_1932_  (.Y(\heichips25_sap3/_1358_ ),
    .A(\heichips25_sap3/sap_3_inst.alu_flags[2] ));
 sg13g2_inv_1 \heichips25_sap3/_1933_  (.Y(\heichips25_sap3/_1359_ ),
    .A(\heichips25_sap3/net1064 ));
 sg13g2_inv_1 \heichips25_sap3/_1934_  (.Y(\heichips25_sap3/_1360_ ),
    .A(\heichips25_sap3/net1130 ));
 sg13g2_inv_1 \heichips25_sap3/_1935_  (.Y(\heichips25_sap3/_1361_ ),
    .A(\heichips25_sap3/net260 ));
 sg13g2_inv_1 \heichips25_sap3/_1936_  (.Y(\heichips25_sap3/_1362_ ),
    .A(\heichips25_sap3/net267 ));
 sg13g2_inv_1 \heichips25_sap3/_1937_  (.Y(\heichips25_sap3/_1363_ ),
    .A(\heichips25_sap3/net264 ));
 sg13g2_inv_1 \heichips25_sap3/_1938_  (.Y(\heichips25_sap3/_1364_ ),
    .A(\heichips25_sap3/net263 ));
 sg13g2_inv_1 \heichips25_sap3/_1939_  (.Y(\heichips25_sap3/_1365_ ),
    .A(\heichips25_sap3/net261 ));
 sg13g2_inv_1 \heichips25_sap3/_1940_  (.Y(\heichips25_sap3/_1366_ ),
    .A(\heichips25_sap3/net830 ));
 sg13g2_inv_1 \heichips25_sap3/_1941_  (.Y(\heichips25_sap3/_1367_ ),
    .A(\heichips25_sap3/net282 ));
 sg13g2_inv_1 \heichips25_sap3/_1942_  (.Y(\heichips25_sap3/_1368_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[0][3] ));
 sg13g2_inv_1 \heichips25_sap3/_1943_  (.Y(\heichips25_sap3/_1369_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][3] ));
 sg13g2_inv_1 \heichips25_sap3/_1944_  (.Y(\heichips25_sap3/_1370_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][3] ));
 sg13g2_inv_1 \heichips25_sap3/_1945_  (.Y(\heichips25_sap3/_1371_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][3] ));
 sg13g2_inv_1 \heichips25_sap3/_1946_  (.Y(\heichips25_sap3/_1372_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][3] ));
 sg13g2_inv_1 \heichips25_sap3/_1947_  (.Y(\heichips25_sap3/_1373_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][3] ));
 sg13g2_inv_1 \heichips25_sap3/_1948_  (.Y(\heichips25_sap3/_1374_ ),
    .A(\heichips25_sap3/net274 ));
 sg13g2_inv_1 \heichips25_sap3/_1949_  (.Y(\heichips25_sap3/_1375_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[0][2] ));
 sg13g2_inv_1 \heichips25_sap3/_1950_  (.Y(\heichips25_sap3/_1376_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][2] ));
 sg13g2_inv_1 \heichips25_sap3/_1951_  (.Y(\heichips25_sap3/_1377_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][2] ));
 sg13g2_inv_1 \heichips25_sap3/_1952_  (.Y(\heichips25_sap3/_1378_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][2] ));
 sg13g2_inv_1 \heichips25_sap3/_1953_  (.Y(\heichips25_sap3/_1379_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][2] ));
 sg13g2_inv_1 \heichips25_sap3/_1954_  (.Y(\heichips25_sap3/_1380_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][2] ));
 sg13g2_inv_1 \heichips25_sap3/_1955_  (.Y(\heichips25_sap3/_1381_ ),
    .A(\heichips25_sap3/net286 ));
 sg13g2_inv_1 \heichips25_sap3/_1956_  (.Y(\heichips25_sap3/_1382_ ),
    .A(\heichips25_sap3/net278 ));
 sg13g2_inv_1 \heichips25_sap3/_1957_  (.Y(\heichips25_sap3/_1383_ ),
    .A(\heichips25_sap3/net280 ));
 sg13g2_inv_1 \heichips25_sap3/_1958_  (.Y(\heichips25_sap3/_1384_ ),
    .A(\heichips25_sap3/net276 ));
 sg13g2_inv_1 \heichips25_sap3/_1959_  (.Y(\heichips25_sap3/_1385_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[0][1] ));
 sg13g2_inv_1 \heichips25_sap3/_1960_  (.Y(\heichips25_sap3/_1386_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][1] ));
 sg13g2_inv_1 \heichips25_sap3/_1961_  (.Y(\heichips25_sap3/_1387_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][1] ));
 sg13g2_inv_1 \heichips25_sap3/_1962_  (.Y(\heichips25_sap3/_1388_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][1] ));
 sg13g2_inv_1 \heichips25_sap3/_1963_  (.Y(\heichips25_sap3/_1389_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][1] ));
 sg13g2_inv_1 \heichips25_sap3/_1964_  (.Y(\heichips25_sap3/_1390_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][1] ));
 sg13g2_inv_1 \heichips25_sap3/_1965_  (.Y(\heichips25_sap3/_1391_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][1] ));
 sg13g2_inv_1 \heichips25_sap3/_1966_  (.Y(\heichips25_sap3/_1392_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[0][0] ));
 sg13g2_inv_1 \heichips25_sap3/_1967_  (.Y(\heichips25_sap3/_1393_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][0] ));
 sg13g2_inv_1 \heichips25_sap3/_1968_  (.Y(\heichips25_sap3/_1394_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][0] ));
 sg13g2_inv_1 \heichips25_sap3/_1969_  (.Y(\heichips25_sap3/_1395_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][0] ));
 sg13g2_inv_1 \heichips25_sap3/_1970_  (.Y(\heichips25_sap3/_1396_ ),
    .A(\heichips25_sap3/sap_3_inst.alu_inst.tmp[1] ));
 sg13g2_inv_1 \heichips25_sap3/_1971_  (.Y(\heichips25_sap3/_1397_ ),
    .A(\heichips25_sap3/sap_3_inst.alu_inst.tmp[2] ));
 sg13g2_inv_1 \heichips25_sap3/_1972_  (.Y(\heichips25_sap3/_1398_ ),
    .A(\heichips25_sap3/sap_3_inst.alu_inst.tmp[6] ));
 sg13g2_inv_1 \heichips25_sap3/_1973_  (.Y(\heichips25_sap3/_1399_ ),
    .A(\heichips25_sap3/sap_3_inst.alu_inst.tmp[7] ));
 sg13g2_inv_1 \heichips25_sap3/_1974_  (.Y(\heichips25_sap3/_1400_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[0][4] ));
 sg13g2_inv_1 \heichips25_sap3/_1975_  (.Y(\heichips25_sap3/_1401_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][4] ));
 sg13g2_inv_1 \heichips25_sap3/_1976_  (.Y(\heichips25_sap3/_1402_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][4] ));
 sg13g2_inv_1 \heichips25_sap3/_1977_  (.Y(\heichips25_sap3/_1403_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][4] ));
 sg13g2_inv_1 \heichips25_sap3/_1978_  (.Y(\heichips25_sap3/_1404_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[0][5] ));
 sg13g2_inv_1 \heichips25_sap3/_1979_  (.Y(\heichips25_sap3/_1405_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][5] ));
 sg13g2_inv_1 \heichips25_sap3/_1980_  (.Y(\heichips25_sap3/_1406_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][5] ));
 sg13g2_inv_1 \heichips25_sap3/_1981_  (.Y(\heichips25_sap3/_1407_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][5] ));
 sg13g2_inv_1 \heichips25_sap3/_1982_  (.Y(\heichips25_sap3/_1408_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][5] ));
 sg13g2_inv_1 \heichips25_sap3/_1983_  (.Y(\heichips25_sap3/_1409_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][5] ));
 sg13g2_inv_1 \heichips25_sap3/_1984_  (.Y(\heichips25_sap3/_1410_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][5] ));
 sg13g2_inv_1 \heichips25_sap3/_1985_  (.Y(\heichips25_sap3/_1411_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][5] ));
 sg13g2_inv_1 \heichips25_sap3/_1986_  (.Y(\heichips25_sap3/_1412_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[0][6] ));
 sg13g2_inv_1 \heichips25_sap3/_1987_  (.Y(\heichips25_sap3/_1413_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][6] ));
 sg13g2_inv_1 \heichips25_sap3/_1988_  (.Y(\heichips25_sap3/_1414_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][6] ));
 sg13g2_inv_1 \heichips25_sap3/_1989_  (.Y(\heichips25_sap3/_1415_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][6] ));
 sg13g2_inv_1 \heichips25_sap3/_1990_  (.Y(\heichips25_sap3/_1416_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][6] ));
 sg13g2_inv_1 \heichips25_sap3/_1991_  (.Y(\heichips25_sap3/_1417_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][6] ));
 sg13g2_inv_1 \heichips25_sap3/_1992_  (.Y(\heichips25_sap3/_1418_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][6] ));
 sg13g2_inv_1 \heichips25_sap3/_1993_  (.Y(\heichips25_sap3/_1419_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][6] ));
 sg13g2_inv_1 \heichips25_sap3/_1994_  (.Y(\heichips25_sap3/_1420_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[0][7] ));
 sg13g2_inv_1 \heichips25_sap3/_1995_  (.Y(\heichips25_sap3/_1421_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][7] ));
 sg13g2_inv_1 \heichips25_sap3/_1996_  (.Y(\heichips25_sap3/_1422_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][7] ));
 sg13g2_inv_1 \heichips25_sap3/_1997_  (.Y(\heichips25_sap3/_1423_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][7] ));
 sg13g2_inv_1 \heichips25_sap3/_1998_  (.Y(\heichips25_sap3/_1424_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][7] ));
 sg13g2_inv_1 \heichips25_sap3/_1999_  (.Y(\heichips25_sap3/_1425_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][7] ));
 sg13g2_inv_1 \heichips25_sap3/_2000_  (.Y(\heichips25_sap3/_1426_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[6] ));
 sg13g2_inv_1 \heichips25_sap3/_2001_  (.Y(\heichips25_sap3/_1427_ ),
    .A(\heichips25_sap3/net1128 ));
 sg13g2_inv_1 \heichips25_sap3/_2002_  (.Y(\heichips25_sap3/_1428_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.word_index[0] ));
 sg13g2_inv_1 \heichips25_sap3/_3871__816  (.Y(net815),
    .A(\clknet_5_25__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_inv_1 \heichips25_sap3/_2004_  (.Y(\heichips25_sap3/_1429_ ),
    .A(\heichips25_sap3/regFile_serial_start ));
 sg13g2_inv_1 \heichips25_sap3/_2005_  (.Y(\heichips25_sap3/_1430_ ),
    .A(\heichips25_sap3/sap_3_outputReg_start_sync ));
 sg13g2_inv_1 \heichips25_sap3/_2006_  (.Y(\heichips25_sap3/u_ser.state[0] ),
    .A(\heichips25_sap3/net341 ));
 sg13g2_inv_1 \heichips25_sap3/_2007_  (.Y(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.state[0] ),
    .A(\heichips25_sap3/net339 ));
 sg13g2_nand2_1 \heichips25_sap3/_2008_  (.Y(\heichips25_sap3/_1431_ ),
    .A(\heichips25_sap3/net1275 ),
    .B(\heichips25_sap3/net1162 ));
 sg13g2_nand2_1 \heichips25_sap3/_2009_  (.Y(\heichips25_sap3/_1432_ ),
    .A(\heichips25_sap3/net1130 ),
    .B(\heichips25_sap3/net835 ));
 sg13g2_or2_1 \heichips25_sap3/_2010_  (.X(\heichips25_sap3/_0018_ ),
    .B(\heichips25_sap3/_1432_ ),
    .A(\heichips25_sap3/_1431_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2011_  (.Y(\heichips25_sap3/_1433_ ),
    .A(\heichips25_sap3/net342 ),
    .B(\heichips25_sap3/net1138 ));
 sg13g2_nand4_1 \heichips25_sap3/_2012_  (.B(\heichips25_sap3/net1019 ),
    .C(\heichips25_sap3/net342 ),
    .A(\heichips25_sap3/u_ser.state[1] ),
    .Y(\heichips25_sap3/_0017_ ),
    .D(\heichips25_sap3/u_ser.bit_pos[1] ));
 sg13g2_nor2_1 \heichips25_sap3/_2013_  (.A(\heichips25_sap3/net258 ),
    .B(\heichips25_sap3/net260 ),
    .Y(\heichips25_sap3/_1434_ ));
 sg13g2_or2_1 \heichips25_sap3/_2014_  (.X(\heichips25_sap3/_1435_ ),
    .B(\heichips25_sap3/net260 ),
    .A(\heichips25_sap3/net258 ));
 sg13g2_nor2_1 \heichips25_sap3/_2015_  (.A(\heichips25_sap3/net267 ),
    .B(\heichips25_sap3/net264 ),
    .Y(\heichips25_sap3/_1436_ ));
 sg13g2_or2_1 \heichips25_sap3/_2016_  (.X(\heichips25_sap3/_1437_ ),
    .B(\heichips25_sap3/net264 ),
    .A(\heichips25_sap3/net267 ));
 sg13g2_or2_1 \heichips25_sap3/_2017_  (.X(\heichips25_sap3/_1438_ ),
    .B(\heichips25_sap3/net261 ),
    .A(\heichips25_sap3/net262 ));
 sg13g2_or2_1 \heichips25_sap3/_2018_  (.X(\heichips25_sap3/_1439_ ),
    .B(\heichips25_sap3/net269 ),
    .A(\heichips25_sap3/net272 ));
 sg13g2_nor4_1 \heichips25_sap3/_2019_  (.A(\heichips25_sap3/_1435_ ),
    .B(\heichips25_sap3/_1437_ ),
    .C(\heichips25_sap3/_1438_ ),
    .D(\heichips25_sap3/_1439_ ),
    .Y(\heichips25_sap3/_1440_ ));
 sg13g2_and2_1 \heichips25_sap3/_2020_  (.A(\heichips25_sap3/net262 ),
    .B(\heichips25_sap3/net261 ),
    .X(\heichips25_sap3/_1441_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2021_  (.Y(\heichips25_sap3/_1442_ ),
    .A(\heichips25_sap3/net263 ),
    .B(\heichips25_sap3/net261 ));
 sg13g2_nor2_1 \heichips25_sap3/_2022_  (.A(\heichips25_sap3/net265 ),
    .B(\heichips25_sap3/net256 ),
    .Y(\heichips25_sap3/_1443_ ));
 sg13g2_nand3b_1 \heichips25_sap3/_2023_  (.B(\heichips25_sap3/net262 ),
    .C(\heichips25_sap3/net261 ),
    .Y(\heichips25_sap3/_1444_ ),
    .A_N(\heichips25_sap3/net264 ));
 sg13g2_nor2b_1 \heichips25_sap3/_2024_  (.A(\heichips25_sap3/net272 ),
    .B_N(\heichips25_sap3/net271 ),
    .Y(\heichips25_sap3/_1445_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_2025_  (.Y(\heichips25_sap3/_1446_ ),
    .B(\heichips25_sap3/net269 ),
    .A_N(\heichips25_sap3/net272 ));
 sg13g2_nor2_1 \heichips25_sap3/_2026_  (.A(\heichips25_sap3/net257 ),
    .B(\heichips25_sap3/_1446_ ),
    .Y(\heichips25_sap3/_1447_ ));
 sg13g2_nand3b_1 \heichips25_sap3/_2027_  (.B(\heichips25_sap3/net269 ),
    .C(\heichips25_sap3/net268 ),
    .Y(\heichips25_sap3/_1448_ ),
    .A_N(\heichips25_sap3/net273 ));
 sg13g2_nor2_1 \heichips25_sap3/_2028_  (.A(\heichips25_sap3/net259 ),
    .B(\heichips25_sap3/_1361_ ),
    .Y(\heichips25_sap3/_1449_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_2029_  (.Y(\heichips25_sap3/_1450_ ),
    .B(\heichips25_sap3/net260 ),
    .A_N(\heichips25_sap3/net259 ));
 sg13g2_nor2_1 \heichips25_sap3/_2030_  (.A(\heichips25_sap3/_1448_ ),
    .B(\heichips25_sap3/_1450_ ),
    .Y(\heichips25_sap3/_1451_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2031_  (.Y(\heichips25_sap3/_1452_ ),
    .A(\heichips25_sap3/_1447_ ),
    .B(\heichips25_sap3/_1449_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2032_  (.A(\heichips25_sap3/_1444_ ),
    .B(\heichips25_sap3/_1450_ ),
    .Y(\heichips25_sap3/_1453_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2033_  (.Y(\heichips25_sap3/_1454_ ),
    .A(\heichips25_sap3/_1443_ ),
    .B(\heichips25_sap3/_1449_ ));
 sg13g2_a21o_1 \heichips25_sap3/_2034_  (.A2(\heichips25_sap3/net248 ),
    .A1(\heichips25_sap3/_1447_ ),
    .B1(\heichips25_sap3/_1440_ ),
    .X(\heichips25_sap3/_1455_ ));
 sg13g2_inv_1 \heichips25_sap3/_2035_  (.Y(\heichips25_sap3/_1456_ ),
    .A(\heichips25_sap3/_1455_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2036_  (.A(\heichips25_sap3/net251 ),
    .B(\heichips25_sap3/net250 ),
    .Y(\heichips25_sap3/_1457_ ));
 sg13g2_or2_1 \heichips25_sap3/_2037_  (.X(\heichips25_sap3/_1458_ ),
    .B(\heichips25_sap3/net250 ),
    .A(\heichips25_sap3/net251 ));
 sg13g2_and2_1 \heichips25_sap3/_2038_  (.A(\heichips25_sap3/net253 ),
    .B(\heichips25_sap3/net252 ),
    .X(\heichips25_sap3/_1459_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2039_  (.Y(\heichips25_sap3/_1460_ ),
    .A(\heichips25_sap3/net253 ),
    .B(\heichips25_sap3/net252 ));
 sg13g2_nor2_1 \heichips25_sap3/_2040_  (.A(\heichips25_sap3/_1458_ ),
    .B(\heichips25_sap3/_1460_ ),
    .Y(\heichips25_sap3/_1461_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2041_  (.Y(\heichips25_sap3/_1462_ ),
    .A(\heichips25_sap3/net247 ),
    .B(\heichips25_sap3/_1459_ ));
 sg13g2_nor2b_1 \heichips25_sap3/_2042_  (.A(\heichips25_sap3/net252 ),
    .B_N(\heichips25_sap3/net253 ),
    .Y(\heichips25_sap3/_1463_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_2043_  (.Y(\heichips25_sap3/_1464_ ),
    .B(\heichips25_sap3/net253 ),
    .A_N(\heichips25_sap3/net252 ));
 sg13g2_nor2_1 \heichips25_sap3/_2044_  (.A(\heichips25_sap3/sap_3_inst.controller_inst.stage[1] ),
    .B(\heichips25_sap3/_1458_ ),
    .Y(\heichips25_sap3/_1465_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2045_  (.Y(\heichips25_sap3/_1466_ ),
    .A(\heichips25_sap3/net247 ),
    .B(\heichips25_sap3/_1463_ ));
 sg13g2_nor2b_1 \heichips25_sap3/_2046_  (.A(\heichips25_sap3/net253 ),
    .B_N(\heichips25_sap3/net252 ),
    .Y(\heichips25_sap3/_1467_ ));
 sg13g2_xor2_1 \heichips25_sap3/_2047_  (.B(\heichips25_sap3/net252 ),
    .A(\heichips25_sap3/net253 ),
    .X(\heichips25_sap3/_1468_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_2048_  (.B2(\heichips25_sap3/net247 ),
    .C1(\heichips25_sap3/_1455_ ),
    .B1(\heichips25_sap3/_1468_ ),
    .A1(\heichips25_sap3/net249 ),
    .Y(\heichips25_sap3/_1469_ ),
    .A2(\heichips25_sap3/net234 ));
 sg13g2_nor2_1 \heichips25_sap3/_2049_  (.A(\heichips25_sap3/_1454_ ),
    .B(\heichips25_sap3/net237 ),
    .Y(\heichips25_sap3/_1470_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_2050_  (.Y(\heichips25_sap3/_1471_ ),
    .B(\heichips25_sap3/_1469_ ),
    .A_N(\heichips25_sap3/_1470_ ));
 sg13g2_nor4_1 \heichips25_sap3/_2051_  (.A(\heichips25_sap3/net257 ),
    .B(\heichips25_sap3/_1435_ ),
    .C(\heichips25_sap3/_1439_ ),
    .D(\heichips25_sap3/_1444_ ),
    .Y(\heichips25_sap3/_1472_ ));
 sg13g2_a21o_1 \heichips25_sap3/_2052_  (.A2(\heichips25_sap3/_1472_ ),
    .A1(\heichips25_sap3/net237 ),
    .B1(\heichips25_sap3/net248 ),
    .X(\heichips25_sap3/_1473_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2053_  (.A(\heichips25_sap3/_1435_ ),
    .B(\heichips25_sap3/_1448_ ),
    .Y(\heichips25_sap3/_1474_ ));
 sg13g2_or2_1 \heichips25_sap3/_2054_  (.X(\heichips25_sap3/_1475_ ),
    .B(\heichips25_sap3/_1448_ ),
    .A(\heichips25_sap3/_1435_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2055_  (.A(\heichips25_sap3/_1444_ ),
    .B(\heichips25_sap3/_1475_ ),
    .Y(\heichips25_sap3/_1476_ ));
 sg13g2_nor2b_1 \heichips25_sap3/_2056_  (.A(\heichips25_sap3/net250 ),
    .B_N(\heichips25_sap3/net251 ),
    .Y(\heichips25_sap3/_1477_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_2057_  (.Y(\heichips25_sap3/_1478_ ),
    .B(\heichips25_sap3/net251 ),
    .A_N(\heichips25_sap3/net250 ));
 sg13g2_nor2_1 \heichips25_sap3/_2058_  (.A(\heichips25_sap3/_1464_ ),
    .B(\heichips25_sap3/_1478_ ),
    .Y(\heichips25_sap3/_1479_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2059_  (.Y(\heichips25_sap3/_1480_ ),
    .A(\heichips25_sap3/_1463_ ),
    .B(\heichips25_sap3/_1477_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2060_  (.Y(\heichips25_sap3/_1481_ ),
    .A(\heichips25_sap3/net234 ),
    .B(\heichips25_sap3/_1480_ ));
 sg13g2_and2_1 \heichips25_sap3/_2061_  (.A(\heichips25_sap3/_1476_ ),
    .B(\heichips25_sap3/_1481_ ),
    .X(\heichips25_sap3/_1482_ ));
 sg13g2_and3_1 \heichips25_sap3/_2062_  (.X(\heichips25_sap3/_1483_ ),
    .A(\heichips25_sap3/net258 ),
    .B(\heichips25_sap3/_1447_ ),
    .C(\heichips25_sap3/net239 ));
 sg13g2_nor3_1 \heichips25_sap3/_2063_  (.A(\heichips25_sap3/_1473_ ),
    .B(\heichips25_sap3/_1482_ ),
    .C(\heichips25_sap3/_1483_ ),
    .Y(\heichips25_sap3/_1484_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2064_  (.A(\heichips25_sap3/_1468_ ),
    .B(\heichips25_sap3/_1478_ ),
    .Y(\heichips25_sap3/_1485_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_2065_  (.Y(\heichips25_sap3/_1486_ ),
    .B(\heichips25_sap3/_1477_ ),
    .A_N(\heichips25_sap3/_1468_ ));
 sg13g2_and2_1 \heichips25_sap3/_2066_  (.A(\heichips25_sap3/net259 ),
    .B(\heichips25_sap3/sap_3_inst.controller_inst.opcode[6] ),
    .X(\heichips25_sap3/_1487_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2067_  (.Y(\heichips25_sap3/_1488_ ),
    .A(\heichips25_sap3/net258 ),
    .B(\heichips25_sap3/net260 ));
 sg13g2_nor2b_1 \heichips25_sap3/_2068_  (.A(\heichips25_sap3/net269 ),
    .B_N(\heichips25_sap3/net273 ),
    .Y(\heichips25_sap3/_1489_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_2069_  (.Y(\heichips25_sap3/_1490_ ),
    .B(\heichips25_sap3/net272 ),
    .A_N(\heichips25_sap3/net271 ));
 sg13g2_nor3_1 \heichips25_sap3/_2070_  (.A(\heichips25_sap3/net257 ),
    .B(\heichips25_sap3/net255 ),
    .C(\heichips25_sap3/_1490_ ),
    .Y(\heichips25_sap3/_1491_ ));
 sg13g2_nand3_1 \heichips25_sap3/_2071_  (.B(\heichips25_sap3/_1487_ ),
    .C(\heichips25_sap3/_1489_ ),
    .A(\heichips25_sap3/net268 ),
    .Y(\heichips25_sap3/_1492_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2072_  (.Y(\heichips25_sap3/_1493_ ),
    .A(\heichips25_sap3/_1485_ ),
    .B(\heichips25_sap3/_1491_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2073_  (.A(\heichips25_sap3/_1437_ ),
    .B(\heichips25_sap3/net255 ),
    .C(\heichips25_sap3/_1490_ ),
    .Y(\heichips25_sap3/_1494_ ));
 sg13g2_nand3_1 \heichips25_sap3/_2074_  (.B(\heichips25_sap3/_1487_ ),
    .C(\heichips25_sap3/_1489_ ),
    .A(\heichips25_sap3/_1436_ ),
    .Y(\heichips25_sap3/_1495_ ));
 sg13g2_and2_1 \heichips25_sap3/_2075_  (.A(\heichips25_sap3/net246 ),
    .B(\heichips25_sap3/_1477_ ),
    .X(\heichips25_sap3/_1496_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2076_  (.Y(\heichips25_sap3/_1497_ ),
    .A(\heichips25_sap3/net246 ),
    .B(\heichips25_sap3/_1477_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2077_  (.A(\heichips25_sap3/net236 ),
    .B(\heichips25_sap3/_1496_ ),
    .Y(\heichips25_sap3/_1498_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2078_  (.Y(\heichips25_sap3/_1499_ ),
    .A(\heichips25_sap3/net235 ),
    .B(\heichips25_sap3/net229 ));
 sg13g2_o21ai_1 \heichips25_sap3/_2079_  (.B1(\heichips25_sap3/_1493_ ),
    .Y(\heichips25_sap3/_1500_ ),
    .A1(\heichips25_sap3/_1495_ ),
    .A2(\heichips25_sap3/_1498_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2080_  (.Y(\heichips25_sap3/_1501_ ),
    .A(\heichips25_sap3/net272 ),
    .B(\heichips25_sap3/net269 ));
 sg13g2_nor2_1 \heichips25_sap3/_2081_  (.A(\heichips25_sap3/_1437_ ),
    .B(\heichips25_sap3/_1501_ ),
    .Y(\heichips25_sap3/_1502_ ));
 sg13g2_nor4_1 \heichips25_sap3/_2082_  (.A(\heichips25_sap3/_1437_ ),
    .B(\heichips25_sap3/_1438_ ),
    .C(\heichips25_sap3/net255 ),
    .D(\heichips25_sap3/_1501_ ),
    .Y(\heichips25_sap3/_1503_ ));
 sg13g2_or4_1 \heichips25_sap3/_2083_  (.A(\heichips25_sap3/_1437_ ),
    .B(\heichips25_sap3/_1438_ ),
    .C(\heichips25_sap3/net255 ),
    .D(\heichips25_sap3/_1501_ ),
    .X(\heichips25_sap3/_1504_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2084_  (.A(\heichips25_sap3/net258 ),
    .B(\heichips25_sap3/net260 ),
    .C(\heichips25_sap3/net267 ),
    .Y(\heichips25_sap3/_1505_ ));
 sg13g2_or3_1 \heichips25_sap3/_2085_  (.A(\heichips25_sap3/net258 ),
    .B(\heichips25_sap3/net260 ),
    .C(\heichips25_sap3/net267 ),
    .X(\heichips25_sap3/_1506_ ));
 sg13g2_nor2b_1 \heichips25_sap3/_2086_  (.A(\heichips25_sap3/net262 ),
    .B_N(\heichips25_sap3/net261 ),
    .Y(\heichips25_sap3/_1507_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_2087_  (.Y(\heichips25_sap3/_1508_ ),
    .B(\heichips25_sap3/net261 ),
    .A_N(\heichips25_sap3/net262 ));
 sg13g2_nor3_1 \heichips25_sap3/_2088_  (.A(\heichips25_sap3/_1446_ ),
    .B(\heichips25_sap3/_1506_ ),
    .C(\heichips25_sap3/_1508_ ),
    .Y(\heichips25_sap3/_1509_ ));
 sg13g2_nand3_1 \heichips25_sap3/_2089_  (.B(\heichips25_sap3/_1505_ ),
    .C(\heichips25_sap3/_1507_ ),
    .A(\heichips25_sap3/_1445_ ),
    .Y(\heichips25_sap3/_1510_ ));
 sg13g2_nand3b_1 \heichips25_sap3/_2090_  (.B(\heichips25_sap3/net266 ),
    .C(\heichips25_sap3/net272 ),
    .Y(\heichips25_sap3/_1511_ ),
    .A_N(\heichips25_sap3/net269 ));
 sg13g2_nor4_2 \heichips25_sap3/_2091_  (.A(\heichips25_sap3/net257 ),
    .B(\heichips25_sap3/_1438_ ),
    .C(\heichips25_sap3/net255 ),
    .Y(\heichips25_sap3/_1512_ ),
    .D(\heichips25_sap3/_1511_ ));
 sg13g2_or4_1 \heichips25_sap3/_2092_  (.A(\heichips25_sap3/net257 ),
    .B(\heichips25_sap3/_1438_ ),
    .C(\heichips25_sap3/net255 ),
    .D(\heichips25_sap3/_1511_ ),
    .X(\heichips25_sap3/_1513_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2093_  (.A(\heichips25_sap3/net245 ),
    .B(\heichips25_sap3/net243 ),
    .Y(\heichips25_sap3/_1514_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2094_  (.A(\heichips25_sap3/net261 ),
    .B(\heichips25_sap3/_1446_ ),
    .C(\heichips25_sap3/_1506_ ),
    .Y(\heichips25_sap3/_1515_ ));
 sg13g2_nand3_1 \heichips25_sap3/_2095_  (.B(\heichips25_sap3/_1445_ ),
    .C(\heichips25_sap3/_1505_ ),
    .A(\heichips25_sap3/_1365_ ),
    .Y(\heichips25_sap3/_1516_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2096_  (.A(\heichips25_sap3/_1506_ ),
    .B(\heichips25_sap3/_1511_ ),
    .Y(\heichips25_sap3/_1517_ ));
 sg13g2_or2_1 \heichips25_sap3/_2097_  (.X(\heichips25_sap3/_1518_ ),
    .B(\heichips25_sap3/_1511_ ),
    .A(\heichips25_sap3/_1506_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2098_  (.A(\heichips25_sap3/_1515_ ),
    .B(\heichips25_sap3/_1517_ ),
    .Y(\heichips25_sap3/_1519_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2099_  (.A(\heichips25_sap3/net256 ),
    .B(\heichips25_sap3/_1446_ ),
    .C(\heichips25_sap3/_1506_ ),
    .Y(\heichips25_sap3/_1520_ ));
 sg13g2_nand3_1 \heichips25_sap3/_2100_  (.B(\heichips25_sap3/_1445_ ),
    .C(\heichips25_sap3/_1505_ ),
    .A(\heichips25_sap3/_1441_ ),
    .Y(\heichips25_sap3/_1521_ ));
 sg13g2_nor4_2 \heichips25_sap3/_2101_  (.A(\heichips25_sap3/net267 ),
    .B(\heichips25_sap3/_1438_ ),
    .C(\heichips25_sap3/_1488_ ),
    .Y(\heichips25_sap3/_1522_ ),
    .D(\heichips25_sap3/_1511_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2102_  (.A(\heichips25_sap3/net242 ),
    .B(\heichips25_sap3/_1522_ ),
    .Y(\heichips25_sap3/_1523_ ));
 sg13g2_and4_1 \heichips25_sap3/_2103_  (.A(\heichips25_sap3/_1504_ ),
    .B(\heichips25_sap3/_1514_ ),
    .C(\heichips25_sap3/_1519_ ),
    .D(\heichips25_sap3/_1523_ ),
    .X(\heichips25_sap3/_1524_ ));
 sg13g2_nand4_1 \heichips25_sap3/_2104_  (.B(\heichips25_sap3/_1514_ ),
    .C(\heichips25_sap3/_1519_ ),
    .A(\heichips25_sap3/_1504_ ),
    .Y(\heichips25_sap3/_1525_ ),
    .D(\heichips25_sap3/_1523_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2105_  (.A(\heichips25_sap3/_1435_ ),
    .B(\heichips25_sap3/_1437_ ),
    .C(\heichips25_sap3/_1490_ ),
    .Y(\heichips25_sap3/_1526_ ));
 sg13g2_nand3_1 \heichips25_sap3/_2106_  (.B(\heichips25_sap3/_1436_ ),
    .C(\heichips25_sap3/_1489_ ),
    .A(\heichips25_sap3/_1434_ ),
    .Y(\heichips25_sap3/_1527_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2107_  (.A(\heichips25_sap3/_1503_ ),
    .B(\heichips25_sap3/_1522_ ),
    .C(\heichips25_sap3/_1526_ ),
    .Y(\heichips25_sap3/_1528_ ));
 sg13g2_nand3b_1 \heichips25_sap3/_2108_  (.B(\heichips25_sap3/net260 ),
    .C(\heichips25_sap3/net258 ),
    .Y(\heichips25_sap3/_1529_ ),
    .A_N(\heichips25_sap3/net272 ));
 sg13g2_nor2_1 \heichips25_sap3/_2109_  (.A(\heichips25_sap3/net267 ),
    .B(\heichips25_sap3/_1529_ ),
    .Y(\heichips25_sap3/_1530_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2110_  (.A(\heichips25_sap3/net257 ),
    .B(\heichips25_sap3/_1439_ ),
    .C(\heichips25_sap3/net255 ),
    .Y(\heichips25_sap3/_1531_ ));
 sg13g2_or3_1 \heichips25_sap3/_2111_  (.A(\heichips25_sap3/net257 ),
    .B(\heichips25_sap3/_1439_ ),
    .C(\heichips25_sap3/net255 ),
    .X(\heichips25_sap3/_1532_ ));
 sg13g2_nor4_1 \heichips25_sap3/_2112_  (.A(\heichips25_sap3/_1474_ ),
    .B(\heichips25_sap3/_1517_ ),
    .C(\heichips25_sap3/_1530_ ),
    .D(\heichips25_sap3/_1531_ ),
    .Y(\heichips25_sap3/_1533_ ));
 sg13g2_and2_1 \heichips25_sap3/_2113_  (.A(\heichips25_sap3/_1528_ ),
    .B(\heichips25_sap3/_1533_ ),
    .X(\heichips25_sap3/_1534_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2114_  (.Y(\heichips25_sap3/_1535_ ),
    .A(\heichips25_sap3/_1528_ ),
    .B(\heichips25_sap3/_1533_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2115_  (.A(\heichips25_sap3/net243 ),
    .B(\heichips25_sap3/_1531_ ),
    .Y(\heichips25_sap3/_1536_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2116_  (.Y(\heichips25_sap3/_1537_ ),
    .A(\heichips25_sap3/_1513_ ),
    .B(\heichips25_sap3/_1532_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2117_  (.A(\heichips25_sap3/_1525_ ),
    .B(\heichips25_sap3/_1535_ ),
    .Y(\heichips25_sap3/_1538_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2118_  (.A(\heichips25_sap3/_1500_ ),
    .B(\heichips25_sap3/_1525_ ),
    .C(\heichips25_sap3/_1535_ ),
    .Y(\heichips25_sap3/_1539_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_2119_  (.Y(\heichips25_sap3/_1540_ ),
    .B(\heichips25_sap3/_1538_ ),
    .A_N(\heichips25_sap3/_1500_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2120_  (.A(\heichips25_sap3/_1364_ ),
    .B(\heichips25_sap3/sap_3_inst.controller_inst.opcode[5] ),
    .Y(\heichips25_sap3/_1541_ ));
 sg13g2_mux4_1 \heichips25_sap3/_2121_  (.S0(\heichips25_sap3/sap_3_inst.controller_inst.opcode[5] ),
    .A0(\heichips25_sap3/sap_3_inst.alu_flags[0] ),
    .A1(\heichips25_sap3/sap_3_inst.alu_flags[2] ),
    .A2(\heichips25_sap3/net254 ),
    .A3(\heichips25_sap3/sap_3_inst.alu_flags[3] ),
    .S1(\heichips25_sap3/net263 ),
    .X(\heichips25_sap3/_1542_ ));
 sg13g2_xnor2_1 \heichips25_sap3/_2122_  (.Y(\heichips25_sap3/_1543_ ),
    .A(\heichips25_sap3/net265 ),
    .B(\heichips25_sap3/_1542_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2123_  (.Y(\heichips25_sap3/_1544_ ),
    .A(\heichips25_sap3/net236 ),
    .B(\heichips25_sap3/_1543_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2124_  (.Y(\heichips25_sap3/_1545_ ),
    .A(\heichips25_sap3/net229 ),
    .B(\heichips25_sap3/_1544_ ));
 sg13g2_nor2b_1 \heichips25_sap3/_2125_  (.A(\heichips25_sap3/net251 ),
    .B_N(\heichips25_sap3/sap_3_inst.controller_inst.stage[3] ),
    .Y(\heichips25_sap3/_1546_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_2126_  (.Y(\heichips25_sap3/_1547_ ),
    .B(\heichips25_sap3/net250 ),
    .A_N(\heichips25_sap3/net251 ));
 sg13g2_nand3b_1 \heichips25_sap3/_2127_  (.B(\heichips25_sap3/sap_3_inst.controller_inst.stage[3] ),
    .C(\heichips25_sap3/net252 ),
    .Y(\heichips25_sap3/_1548_ ),
    .A_N(\heichips25_sap3/sap_3_inst.controller_inst.stage[2] ));
 sg13g2_nor2_1 \heichips25_sap3/_2128_  (.A(\heichips25_sap3/net253 ),
    .B(\heichips25_sap3/_1548_ ),
    .Y(\heichips25_sap3/_1549_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2129_  (.Y(\heichips25_sap3/_1550_ ),
    .A(\heichips25_sap3/net246 ),
    .B(\heichips25_sap3/_1546_ ));
 sg13g2_and2_1 \heichips25_sap3/_2130_  (.A(\heichips25_sap3/net251 ),
    .B(\heichips25_sap3/net250 ),
    .X(\heichips25_sap3/_1551_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2131_  (.Y(\heichips25_sap3/_1552_ ),
    .A(\heichips25_sap3/net251 ),
    .B(\heichips25_sap3/net250 ));
 sg13g2_a22oi_1 \heichips25_sap3/_2132_  (.Y(\heichips25_sap3/_1553_ ),
    .B1(\heichips25_sap3/_1551_ ),
    .B2(\heichips25_sap3/_1463_ ),
    .A2(\heichips25_sap3/_1546_ ),
    .A1(\heichips25_sap3/net246 ));
 sg13g2_nand2_1 \heichips25_sap3/_2133_  (.Y(\heichips25_sap3/_1554_ ),
    .A(\heichips25_sap3/sap_3_inst.controller_inst.stage[2] ),
    .B(\heichips25_sap3/_1459_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2134_  (.B1(\heichips25_sap3/_1553_ ),
    .Y(\heichips25_sap3/_1555_ ),
    .A1(\heichips25_sap3/_1460_ ),
    .A2(\heichips25_sap3/_1552_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2135_  (.B1(\heichips25_sap3/_1531_ ),
    .Y(\heichips25_sap3/_1556_ ),
    .A1(\heichips25_sap3/_1545_ ),
    .A2(\heichips25_sap3/_1555_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2136_  (.A(\heichips25_sap3/net267 ),
    .B(\heichips25_sap3/net269 ),
    .C(\heichips25_sap3/_1529_ ),
    .Y(\heichips25_sap3/_1557_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_2137_  (.Y(\heichips25_sap3/_1558_ ),
    .B(\heichips25_sap3/_1530_ ),
    .A_N(\heichips25_sap3/net271 ));
 sg13g2_nor2_1 \heichips25_sap3/_2138_  (.A(\heichips25_sap3/_1464_ ),
    .B(\heichips25_sap3/_1547_ ),
    .Y(\heichips25_sap3/_1559_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2139_  (.Y(\heichips25_sap3/_1560_ ),
    .A(\heichips25_sap3/_1463_ ),
    .B(\heichips25_sap3/_1546_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2140_  (.A(\heichips25_sap3/_1496_ ),
    .B(\heichips25_sap3/_1559_ ),
    .Y(\heichips25_sap3/_1561_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2141_  (.A1(\heichips25_sap3/_1544_ ),
    .A2(\heichips25_sap3/_1561_ ),
    .Y(\heichips25_sap3/_1562_ ),
    .B1(\heichips25_sap3/_1558_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2142_  (.Y(\heichips25_sap3/_1563_ ),
    .A(\heichips25_sap3/_1498_ ),
    .B(\heichips25_sap3/_1560_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_2143_  (.B2(\heichips25_sap3/_1522_ ),
    .C1(\heichips25_sap3/_1562_ ),
    .B1(\heichips25_sap3/_1563_ ),
    .A1(\heichips25_sap3/_1524_ ),
    .Y(\heichips25_sap3/_1564_ ),
    .A2(\heichips25_sap3/_1534_ ));
 sg13g2_nand3b_1 \heichips25_sap3/_2144_  (.B(\heichips25_sap3/net257 ),
    .C(\heichips25_sap3/net269 ),
    .Y(\heichips25_sap3/_1565_ ),
    .A_N(\heichips25_sap3/_1529_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2145_  (.A(\heichips25_sap3/sap_3_inst.controller_inst.stage[0] ),
    .B(\heichips25_sap3/sap_3_inst.controller_inst.stage[1] ),
    .Y(\heichips25_sap3/_1566_ ));
 sg13g2_or2_1 \heichips25_sap3/_2146_  (.X(\heichips25_sap3/_1567_ ),
    .B(\heichips25_sap3/net252 ),
    .A(\heichips25_sap3/net253 ));
 sg13g2_nor2_1 \heichips25_sap3/_2147_  (.A(\heichips25_sap3/_1547_ ),
    .B(\heichips25_sap3/_1567_ ),
    .Y(\heichips25_sap3/_1568_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2148_  (.Y(\heichips25_sap3/_1569_ ),
    .A(\heichips25_sap3/_1546_ ),
    .B(\heichips25_sap3/_1566_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2149_  (.A(\heichips25_sap3/_1496_ ),
    .B(\heichips25_sap3/_1568_ ),
    .Y(\heichips25_sap3/_1570_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2150_  (.A1(\heichips25_sap3/_1544_ ),
    .A2(\heichips25_sap3/_1570_ ),
    .Y(\heichips25_sap3/_1571_ ),
    .B1(\heichips25_sap3/_1565_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2151_  (.Y(\heichips25_sap3/_1572_ ),
    .A(\heichips25_sap3/_1459_ ),
    .B(\heichips25_sap3/_1546_ ));
 sg13g2_or4_1 \heichips25_sap3/_2152_  (.A(\heichips25_sap3/_1460_ ),
    .B(\heichips25_sap3/_1506_ ),
    .C(\heichips25_sap3/_1511_ ),
    .D(\heichips25_sap3/_1547_ ),
    .X(\heichips25_sap3/_1573_ ));
 sg13g2_inv_1 \heichips25_sap3/_2153_  (.Y(\heichips25_sap3/_1574_ ),
    .A(\heichips25_sap3/_1573_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2154_  (.A1(\heichips25_sap3/net229 ),
    .A2(\heichips25_sap3/_1553_ ),
    .Y(\heichips25_sap3/_1575_ ),
    .B1(\heichips25_sap3/_1513_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2155_  (.A1(\heichips25_sap3/_1458_ ),
    .A2(\heichips25_sap3/_1552_ ),
    .Y(\heichips25_sap3/_1576_ ),
    .B1(\heichips25_sap3/_1460_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2156_  (.A(\heichips25_sap3/_1480_ ),
    .B(\heichips25_sap3/_1516_ ),
    .Y(\heichips25_sap3/_1577_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2157_  (.A(\heichips25_sap3/net234 ),
    .B(\heichips25_sap3/_1475_ ),
    .Y(\heichips25_sap3/_1578_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2158_  (.A(\heichips25_sap3/_1577_ ),
    .B(\heichips25_sap3/_1578_ ),
    .Y(\heichips25_sap3/_1579_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2159_  (.Y(\heichips25_sap3/_1580_ ),
    .B1(\heichips25_sap3/_1551_ ),
    .B2(\heichips25_sap3/_1566_ ),
    .A2(\heichips25_sap3/_1546_ ),
    .A1(\heichips25_sap3/_1463_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2160_  (.B1(\heichips25_sap3/_1560_ ),
    .Y(\heichips25_sap3/_1581_ ),
    .A1(\heichips25_sap3/_1552_ ),
    .A2(\heichips25_sap3/_1567_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2161_  (.B1(\heichips25_sap3/net245 ),
    .Y(\heichips25_sap3/_1582_ ),
    .A1(\heichips25_sap3/_1499_ ),
    .A2(\heichips25_sap3/_1581_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2162_  (.Y(\heichips25_sap3/_1583_ ),
    .B1(\heichips25_sap3/_1569_ ),
    .B2(\heichips25_sap3/_1498_ ),
    .A2(\heichips25_sap3/_1527_ ),
    .A1(\heichips25_sap3/_1504_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_2163_  (.Y(\heichips25_sap3/_1584_ ),
    .B(\heichips25_sap3/_1582_ ),
    .A_N(\heichips25_sap3/_1575_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2164_  (.Y(\heichips25_sap3/_1585_ ),
    .B1(\heichips25_sap3/_1576_ ),
    .B2(\heichips25_sap3/net243 ),
    .A2(\heichips25_sap3/_1563_ ),
    .A1(\heichips25_sap3/net242 ));
 sg13g2_nor2_1 \heichips25_sap3/_2165_  (.A(\heichips25_sap3/_1574_ ),
    .B(\heichips25_sap3/_1583_ ),
    .Y(\heichips25_sap3/_1586_ ));
 sg13g2_nand3_1 \heichips25_sap3/_2166_  (.B(\heichips25_sap3/_1585_ ),
    .C(\heichips25_sap3/_1586_ ),
    .A(\heichips25_sap3/_1579_ ),
    .Y(\heichips25_sap3/_1587_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2167_  (.A(\heichips25_sap3/_1571_ ),
    .B(\heichips25_sap3/_1584_ ),
    .C(\heichips25_sap3/_1587_ ),
    .Y(\heichips25_sap3/_1588_ ));
 sg13g2_nand3_1 \heichips25_sap3/_2168_  (.B(\heichips25_sap3/_1564_ ),
    .C(\heichips25_sap3/_1588_ ),
    .A(\heichips25_sap3/_1556_ ),
    .Y(\heichips25_sap3/_1589_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2169_  (.Y(\heichips25_sap3/_1590_ ),
    .A(\heichips25_sap3/_1540_ ),
    .B(\heichips25_sap3/_1589_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2170_  (.A1(\heichips25_sap3/_1484_ ),
    .A2(\heichips25_sap3/_1590_ ),
    .Y(\heichips25_sap3/_1591_ ),
    .B1(\heichips25_sap3/_1471_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2171_  (.Y(\heichips25_sap3/_1592_ ),
    .A(\heichips25_sap3/net247 ),
    .B(\heichips25_sap3/_1566_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_2172_  (.B2(\heichips25_sap3/net247 ),
    .C1(\heichips25_sap3/_1591_ ),
    .B1(\heichips25_sap3/_1566_ ),
    .A1(\heichips25_sap3/net249 ),
    .Y(\heichips25_sap3/_1593_ ),
    .A2(\heichips25_sap3/_1469_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2173_  (.B1(\heichips25_sap3/_1526_ ),
    .Y(\heichips25_sap3/_1594_ ),
    .A1(\heichips25_sap3/_1499_ ),
    .A2(\heichips25_sap3/_1568_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2174_  (.A1(\heichips25_sap3/_1504_ ),
    .A2(\heichips25_sap3/_1525_ ),
    .Y(\heichips25_sap3/_1595_ ),
    .B1(\heichips25_sap3/_1570_ ));
 sg13g2_inv_1 \heichips25_sap3/_2175_  (.Y(\heichips25_sap3/_1596_ ),
    .A(\heichips25_sap3/_1595_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2176_  (.A(\heichips25_sap3/_1478_ ),
    .B(\heichips25_sap3/_1567_ ),
    .Y(\heichips25_sap3/_1597_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2177_  (.Y(\heichips25_sap3/_1598_ ),
    .A(\heichips25_sap3/_1477_ ),
    .B(\heichips25_sap3/_1566_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2178_  (.A(\heichips25_sap3/_1519_ ),
    .B(\heichips25_sap3/net225 ),
    .Y(\heichips25_sap3/_1599_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2179_  (.A(\heichips25_sap3/_1523_ ),
    .B(\heichips25_sap3/_1561_ ),
    .Y(\heichips25_sap3/_1600_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2180_  (.A(\heichips25_sap3/net266 ),
    .B(\heichips25_sap3/_1510_ ),
    .C(\heichips25_sap3/_1553_ ),
    .Y(\heichips25_sap3/_1601_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2181_  (.Y(\heichips25_sap3/_1602_ ),
    .A(\heichips25_sap3/_1551_ ),
    .B(\heichips25_sap3/_1567_ ));
 sg13g2_nand3_1 \heichips25_sap3/_2182_  (.B(\heichips25_sap3/_1548_ ),
    .C(\heichips25_sap3/_1602_ ),
    .A(\heichips25_sap3/net229 ),
    .Y(\heichips25_sap3/_1603_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2183_  (.A1(\heichips25_sap3/net243 ),
    .A2(\heichips25_sap3/_1603_ ),
    .Y(\heichips25_sap3/_1604_ ),
    .B1(\heichips25_sap3/_1577_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2184_  (.A(\heichips25_sap3/_1460_ ),
    .B(\heichips25_sap3/_1478_ ),
    .Y(\heichips25_sap3/_1605_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2185_  (.Y(\heichips25_sap3/_1606_ ),
    .A(\heichips25_sap3/_1459_ ),
    .B(\heichips25_sap3/_1477_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2186_  (.A(\heichips25_sap3/_1468_ ),
    .B(\heichips25_sap3/_1547_ ),
    .Y(\heichips25_sap3/_1607_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2187_  (.B1(\heichips25_sap3/_1517_ ),
    .Y(\heichips25_sap3/_1608_ ),
    .A1(\heichips25_sap3/_1605_ ),
    .A2(\heichips25_sap3/_1607_ ));
 sg13g2_nand4_1 \heichips25_sap3/_2188_  (.B(\heichips25_sap3/_1582_ ),
    .C(\heichips25_sap3/_1604_ ),
    .A(\heichips25_sap3/net235 ),
    .Y(\heichips25_sap3/_1609_ ),
    .D(\heichips25_sap3/_1608_ ));
 sg13g2_nor4_1 \heichips25_sap3/_2189_  (.A(\heichips25_sap3/_1599_ ),
    .B(\heichips25_sap3/_1600_ ),
    .C(\heichips25_sap3/_1601_ ),
    .D(\heichips25_sap3/_1609_ ),
    .Y(\heichips25_sap3/_1610_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2190_  (.Y(\heichips25_sap3/_1611_ ),
    .B1(\heichips25_sap3/_1596_ ),
    .B2(\heichips25_sap3/_1610_ ),
    .A2(\heichips25_sap3/_1594_ ),
    .A1(\heichips25_sap3/_1524_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2191_  (.Y(\heichips25_sap3/_1612_ ),
    .A(\heichips25_sap3/_1500_ ),
    .B(\heichips25_sap3/_1513_ ));
 sg13g2_nand3_1 \heichips25_sap3/_2192_  (.B(\heichips25_sap3/net273 ),
    .C(\heichips25_sap3/net270 ),
    .A(\heichips25_sap3/net268 ),
    .Y(\heichips25_sap3/_1613_ ));
 sg13g2_nor2b_1 \heichips25_sap3/_2193_  (.A(\heichips25_sap3/sap_3_inst.controller_inst.opcode[6] ),
    .B_N(\heichips25_sap3/net259 ),
    .Y(\heichips25_sap3/_1614_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_2194_  (.Y(\heichips25_sap3/_1615_ ),
    .B(\heichips25_sap3/net259 ),
    .A_N(\heichips25_sap3/sap_3_inst.controller_inst.opcode[6] ));
 sg13g2_nand2_1 \heichips25_sap3/_2195_  (.Y(\heichips25_sap3/_1616_ ),
    .A(\heichips25_sap3/net237 ),
    .B(\heichips25_sap3/_1613_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2196_  (.A(\heichips25_sap3/_1615_ ),
    .B(\heichips25_sap3/_1616_ ),
    .Y(\heichips25_sap3/_1617_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2197_  (.A(\heichips25_sap3/_1362_ ),
    .B(\heichips25_sap3/net270 ),
    .C(\heichips25_sap3/_1435_ ),
    .Y(\heichips25_sap3/_1618_ ));
 sg13g2_nand3b_1 \heichips25_sap3/_2198_  (.B(\heichips25_sap3/_1434_ ),
    .C(\heichips25_sap3/net268 ),
    .Y(\heichips25_sap3/_1619_ ),
    .A_N(\heichips25_sap3/net270 ));
 sg13g2_nor2_1 \heichips25_sap3/_2199_  (.A(\heichips25_sap3/_1448_ ),
    .B(\heichips25_sap3/_1615_ ),
    .Y(\heichips25_sap3/_1620_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2200_  (.A(\heichips25_sap3/_1618_ ),
    .B(\heichips25_sap3/_1620_ ),
    .Y(\heichips25_sap3/_1621_ ));
 sg13g2_or2_1 \heichips25_sap3/_2201_  (.X(\heichips25_sap3/_1622_ ),
    .B(\heichips25_sap3/_1620_ ),
    .A(\heichips25_sap3/_1618_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2202_  (.A(\heichips25_sap3/_1448_ ),
    .B(\heichips25_sap3/_1488_ ),
    .Y(\heichips25_sap3/_1623_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2203_  (.Y(\heichips25_sap3/_1624_ ),
    .A(\heichips25_sap3/net240 ),
    .B(\heichips25_sap3/_1623_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2204_  (.Y(\heichips25_sap3/_1625_ ),
    .B1(\heichips25_sap3/_1546_ ),
    .B2(\heichips25_sap3/_1566_ ),
    .A2(\heichips25_sap3/_1477_ ),
    .A1(\heichips25_sap3/_1463_ ));
 sg13g2_inv_1 \heichips25_sap3/_2205_  (.Y(\heichips25_sap3/_1626_ ),
    .A(\heichips25_sap3/net222 ));
 sg13g2_nor2_1 \heichips25_sap3/_2206_  (.A(\heichips25_sap3/_1492_ ),
    .B(\heichips25_sap3/net222 ),
    .Y(\heichips25_sap3/_1627_ ));
 sg13g2_nor4_1 \heichips25_sap3/_2207_  (.A(\heichips25_sap3/_1441_ ),
    .B(\heichips25_sap3/_1492_ ),
    .C(\heichips25_sap3/net244 ),
    .D(\heichips25_sap3/net222 ),
    .Y(\heichips25_sap3/_1628_ ));
 sg13g2_nand3_1 \heichips25_sap3/_2208_  (.B(\heichips25_sap3/_1476_ ),
    .C(\heichips25_sap3/_1477_ ),
    .A(\heichips25_sap3/net246 ),
    .Y(\heichips25_sap3/_1629_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2209_  (.Y(\heichips25_sap3/_1630_ ),
    .A(\heichips25_sap3/_1476_ ),
    .B(\heichips25_sap3/_1496_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2210_  (.A(\heichips25_sap3/_1482_ ),
    .B(\heichips25_sap3/net223 ),
    .Y(\heichips25_sap3/_1631_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2211_  (.A(\heichips25_sap3/_1448_ ),
    .B(\heichips25_sap3/net234 ),
    .C(\heichips25_sap3/_1488_ ),
    .Y(\heichips25_sap3/_1632_ ));
 sg13g2_nor4_1 \heichips25_sap3/_2212_  (.A(\heichips25_sap3/_1578_ ),
    .B(\heichips25_sap3/_1617_ ),
    .C(\heichips25_sap3/_1628_ ),
    .D(\heichips25_sap3/_1632_ ),
    .Y(\heichips25_sap3/_1633_ ));
 sg13g2_nand4_1 \heichips25_sap3/_2213_  (.B(\heichips25_sap3/_1630_ ),
    .C(\heichips25_sap3/_1631_ ),
    .A(\heichips25_sap3/_1612_ ),
    .Y(\heichips25_sap3/_1634_ ),
    .D(\heichips25_sap3/_1633_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_2214_  (.Y(\heichips25_sap3/_1635_ ),
    .B(\heichips25_sap3/net236 ),
    .A_N(\heichips25_sap3/_1543_ ));
 sg13g2_and2_1 \heichips25_sap3/_2215_  (.A(\heichips25_sap3/_1531_ ),
    .B(\heichips25_sap3/_1635_ ),
    .X(\heichips25_sap3/_1636_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2216_  (.B1(\heichips25_sap3/_1636_ ),
    .Y(\heichips25_sap3/_1637_ ),
    .A1(\heichips25_sap3/net236 ),
    .A2(\heichips25_sap3/_1603_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_2217_  (.Y(\heichips25_sap3/_1638_ ),
    .B(\heichips25_sap3/_1637_ ),
    .A_N(\heichips25_sap3/_1571_ ));
 sg13g2_nor4_1 \heichips25_sap3/_2218_  (.A(\heichips25_sap3/_1562_ ),
    .B(\heichips25_sap3/_1611_ ),
    .C(\heichips25_sap3/_1634_ ),
    .D(\heichips25_sap3/_1638_ ),
    .Y(\heichips25_sap3/_1639_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2219_  (.B1(\heichips25_sap3/_1450_ ),
    .Y(\heichips25_sap3/_1640_ ),
    .A1(\heichips25_sap3/_1501_ ),
    .A2(\heichips25_sap3/_1506_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2220_  (.A(\heichips25_sap3/_1472_ ),
    .B(\heichips25_sap3/_1640_ ),
    .Y(\heichips25_sap3/_1641_ ));
 sg13g2_or2_1 \heichips25_sap3/_2221_  (.X(\heichips25_sap3/_1642_ ),
    .B(\heichips25_sap3/_1640_ ),
    .A(\heichips25_sap3/_1472_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2222_  (.A(\heichips25_sap3/_1363_ ),
    .B(\heichips25_sap3/net256 ),
    .Y(\heichips25_sap3/_1643_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2223_  (.Y(\heichips25_sap3/_1644_ ),
    .A(\heichips25_sap3/net264 ),
    .B(\heichips25_sap3/_1441_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2224_  (.Y(\heichips25_sap3/_1645_ ),
    .A(\heichips25_sap3/net238 ),
    .B(\heichips25_sap3/_1644_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2225_  (.B1(\heichips25_sap3/net223 ),
    .Y(\heichips25_sap3/_1646_ ),
    .A1(\heichips25_sap3/_1619_ ),
    .A2(\heichips25_sap3/_1645_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2226_  (.A1(\heichips25_sap3/net237 ),
    .A2(\heichips25_sap3/_1620_ ),
    .Y(\heichips25_sap3/_1647_ ),
    .B1(\heichips25_sap3/_1646_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2227_  (.A(\heichips25_sap3/_1639_ ),
    .B(\heichips25_sap3/net220 ),
    .C(\heichips25_sap3/_1647_ ),
    .Y(\heichips25_sap3/_1648_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2228_  (.A(\heichips25_sap3/_1450_ ),
    .B(\heichips25_sap3/_1616_ ),
    .Y(\heichips25_sap3/_1649_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2229_  (.A(\heichips25_sap3/_1473_ ),
    .B(\heichips25_sap3/_1648_ ),
    .C(\heichips25_sap3/_1649_ ),
    .Y(\heichips25_sap3/_1650_ ));
 sg13g2_and2_1 \heichips25_sap3/_2230_  (.A(\heichips25_sap3/net227 ),
    .B(\heichips25_sap3/_1613_ ),
    .X(\heichips25_sap3/_1651_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2231_  (.Y(\heichips25_sap3/_1652_ ),
    .A(\heichips25_sap3/_1469_ ),
    .B(\heichips25_sap3/_1651_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2232_  (.Y(\heichips25_sap3/_1653_ ),
    .A(\heichips25_sap3/_1471_ ),
    .B(\heichips25_sap3/_1652_ ));
 sg13g2_nand3b_1 \heichips25_sap3/_2233_  (.B(\heichips25_sap3/_1653_ ),
    .C(\heichips25_sap3/net67 ),
    .Y(\heichips25_sap3/_1654_ ),
    .A_N(\heichips25_sap3/_1650_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2234_  (.Y(\heichips25_sap3/_1655_ ),
    .A(\heichips25_sap3/net268 ),
    .B(\heichips25_sap3/_1501_ ));
 sg13g2_inv_1 \heichips25_sap3/_2235_  (.Y(\heichips25_sap3/_1656_ ),
    .A(\heichips25_sap3/_1655_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2236_  (.A1(\heichips25_sap3/net238 ),
    .A2(\heichips25_sap3/_1656_ ),
    .Y(\heichips25_sap3/_1657_ ),
    .B1(\heichips25_sap3/_1641_ ));
 sg13g2_nand3_1 \heichips25_sap3/_2237_  (.B(\heichips25_sap3/_1527_ ),
    .C(\heichips25_sap3/_1565_ ),
    .A(\heichips25_sap3/_1504_ ),
    .Y(\heichips25_sap3/_1658_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2238_  (.Y(\heichips25_sap3/_1659_ ),
    .A(\heichips25_sap3/_1568_ ),
    .B(\heichips25_sap3/_1658_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_2239_  (.B2(\heichips25_sap3/net245 ),
    .C1(\heichips25_sap3/_1577_ ),
    .B1(\heichips25_sap3/_1581_ ),
    .A1(\heichips25_sap3/net242 ),
    .Y(\heichips25_sap3/_1660_ ),
    .A2(\heichips25_sap3/_1559_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2240_  (.Y(\heichips25_sap3/_1661_ ),
    .A(\heichips25_sap3/_1659_ ),
    .B(\heichips25_sap3/_1660_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2241_  (.A1(\heichips25_sap3/_1569_ ),
    .A2(\heichips25_sap3/net225 ),
    .Y(\heichips25_sap3/_1662_ ),
    .B1(\heichips25_sap3/_1518_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2242_  (.B1(\heichips25_sap3/_1507_ ),
    .Y(\heichips25_sap3/_1663_ ),
    .A1(\heichips25_sap3/_1627_ ),
    .A2(\heichips25_sap3/_1662_ ));
 sg13g2_or2_1 \heichips25_sap3/_2243_  (.X(\heichips25_sap3/_1664_ ),
    .B(\heichips25_sap3/_1557_ ),
    .A(\heichips25_sap3/_1522_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2244_  (.Y(\heichips25_sap3/_1665_ ),
    .A(\heichips25_sap3/_1559_ ),
    .B(\heichips25_sap3/_1664_ ));
 sg13g2_nand3_1 \heichips25_sap3/_2245_  (.B(\heichips25_sap3/_1537_ ),
    .C(\heichips25_sap3/_1551_ ),
    .A(\heichips25_sap3/_1459_ ),
    .Y(\heichips25_sap3/_1666_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2246_  (.A(\heichips25_sap3/_1601_ ),
    .B(\heichips25_sap3/net220 ),
    .Y(\heichips25_sap3/_1667_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2247_  (.A1(\heichips25_sap3/net266 ),
    .A2(\heichips25_sap3/net262 ),
    .Y(\heichips25_sap3/_1668_ ),
    .B1(\heichips25_sap3/_1365_ ));
 sg13g2_nand3_1 \heichips25_sap3/_2248_  (.B(\heichips25_sap3/net223 ),
    .C(\heichips25_sap3/_1668_ ),
    .A(\heichips25_sap3/net240 ),
    .Y(\heichips25_sap3/_1669_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2249_  (.A(\heichips25_sap3/net250 ),
    .B(\heichips25_sap3/_1460_ ),
    .C(\heichips25_sap3/_1518_ ),
    .Y(\heichips25_sap3/_1670_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2250_  (.A(\heichips25_sap3/_1462_ ),
    .B(\heichips25_sap3/_1615_ ),
    .C(\heichips25_sap3/_1655_ ),
    .Y(\heichips25_sap3/_1671_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2251_  (.A(\heichips25_sap3/_1574_ ),
    .B(\heichips25_sap3/_1670_ ),
    .C(\heichips25_sap3/_1671_ ),
    .Y(\heichips25_sap3/_1672_ ));
 sg13g2_nand4_1 \heichips25_sap3/_2252_  (.B(\heichips25_sap3/_1666_ ),
    .C(\heichips25_sap3/_1669_ ),
    .A(\heichips25_sap3/_1663_ ),
    .Y(\heichips25_sap3/_1673_ ),
    .D(\heichips25_sap3/_1672_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2253_  (.B1(\heichips25_sap3/_1476_ ),
    .Y(\heichips25_sap3/_1674_ ),
    .A1(\heichips25_sap3/net230 ),
    .A2(\heichips25_sap3/_1496_ ));
 sg13g2_nand3_1 \heichips25_sap3/_2254_  (.B(\heichips25_sap3/_1667_ ),
    .C(\heichips25_sap3/_1674_ ),
    .A(\heichips25_sap3/_1665_ ),
    .Y(\heichips25_sap3/_1675_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2255_  (.A(\heichips25_sap3/_1661_ ),
    .B(\heichips25_sap3/_1673_ ),
    .C(\heichips25_sap3/_1675_ ),
    .Y(\heichips25_sap3/_1676_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2256_  (.B1(\heichips25_sap3/_1454_ ),
    .Y(\heichips25_sap3/_1677_ ),
    .A1(\heichips25_sap3/_1657_ ),
    .A2(\heichips25_sap3/_1676_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2257_  (.B1(\heichips25_sap3/_1470_ ),
    .Y(\heichips25_sap3/_1678_ ),
    .A1(\heichips25_sap3/net225 ),
    .A2(\heichips25_sap3/_1655_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2258_  (.Y(\heichips25_sap3/_1679_ ),
    .A(\heichips25_sap3/net247 ),
    .B(\heichips25_sap3/_1460_ ));
 sg13g2_and4_1 \heichips25_sap3/_2259_  (.A(\heichips25_sap3/_1456_ ),
    .B(\heichips25_sap3/_1677_ ),
    .C(\heichips25_sap3/_1678_ ),
    .D(\heichips25_sap3/_1679_ ),
    .X(\heichips25_sap3/_1680_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2260_  (.Y(\heichips25_sap3/_1681_ ),
    .B1(\heichips25_sap3/_1551_ ),
    .B2(\heichips25_sap3/net246 ),
    .A2(\heichips25_sap3/_1546_ ),
    .A1(\heichips25_sap3/_1459_ ));
 sg13g2_inv_1 \heichips25_sap3/_2261_  (.Y(\heichips25_sap3/_1682_ ),
    .A(\heichips25_sap3/_1681_ ));
 sg13g2_nand4_1 \heichips25_sap3/_2262_  (.B(\heichips25_sap3/_1544_ ),
    .C(\heichips25_sap3/_1553_ ),
    .A(\heichips25_sap3/net229 ),
    .Y(\heichips25_sap3/_1683_ ),
    .D(\heichips25_sap3/_1681_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2263_  (.Y(\heichips25_sap3/_1684_ ),
    .B1(\heichips25_sap3/_1683_ ),
    .B2(\heichips25_sap3/_1531_ ),
    .A2(\heichips25_sap3/_1545_ ),
    .A1(\heichips25_sap3/_1530_ ));
 sg13g2_nor4_1 \heichips25_sap3/_2264_  (.A(\heichips25_sap3/_1503_ ),
    .B(\heichips25_sap3/net242 ),
    .C(\heichips25_sap3/_1522_ ),
    .D(\heichips25_sap3/_1526_ ),
    .Y(\heichips25_sap3/_1685_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2265_  (.A1(\heichips25_sap3/net236 ),
    .A2(\heichips25_sap3/_1474_ ),
    .Y(\heichips25_sap3/_1686_ ),
    .B1(\heichips25_sap3/net245 ));
 sg13g2_nand2_1 \heichips25_sap3/_2266_  (.Y(\heichips25_sap3/_1687_ ),
    .A(\heichips25_sap3/_1685_ ),
    .B(\heichips25_sap3/_1686_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2267_  (.Y(\heichips25_sap3/_1688_ ),
    .A(\heichips25_sap3/_1441_ ),
    .B(\heichips25_sap3/_1662_ ));
 sg13g2_nand4_1 \heichips25_sap3/_2268_  (.B(\heichips25_sap3/net229 ),
    .C(\heichips25_sap3/_1553_ ),
    .A(\heichips25_sap3/net235 ),
    .Y(\heichips25_sap3/_1689_ ),
    .D(\heichips25_sap3/_1681_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2269_  (.Y(\heichips25_sap3/_1690_ ),
    .B1(\heichips25_sap3/_1689_ ),
    .B2(\heichips25_sap3/net243 ),
    .A2(\heichips25_sap3/_1687_ ),
    .A1(\heichips25_sap3/_1499_ ));
 sg13g2_nand3_1 \heichips25_sap3/_2270_  (.B(\heichips25_sap3/_1688_ ),
    .C(\heichips25_sap3/_1690_ ),
    .A(\heichips25_sap3/_1684_ ),
    .Y(\heichips25_sap3/_1691_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2271_  (.B1(\heichips25_sap3/_1540_ ),
    .Y(\heichips25_sap3/_1692_ ),
    .A1(\heichips25_sap3/_1538_ ),
    .A2(\heichips25_sap3/_1691_ ));
 sg13g2_nand3_1 \heichips25_sap3/_2272_  (.B(\heichips25_sap3/_1624_ ),
    .C(\heichips25_sap3/_1692_ ),
    .A(\heichips25_sap3/_1592_ ),
    .Y(\heichips25_sap3/_1693_ ));
 sg13g2_inv_1 \heichips25_sap3/_2273_  (.Y(\heichips25_sap3/_1694_ ),
    .A(\heichips25_sap3/_1693_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2274_  (.A(\heichips25_sap3/_1680_ ),
    .B(\heichips25_sap3/_1693_ ),
    .Y(\heichips25_sap3/_1695_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2275_  (.Y(\heichips25_sap3/_1696_ ),
    .A(\heichips25_sap3/_1541_ ),
    .B(\heichips25_sap3/_1627_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2276_  (.A1(\heichips25_sap3/net234 ),
    .A2(\heichips25_sap3/net225 ),
    .Y(\heichips25_sap3/_1697_ ),
    .B1(\heichips25_sap3/_1516_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2277_  (.B1(\heichips25_sap3/_1697_ ),
    .Y(\heichips25_sap3/_1698_ ),
    .A1(\heichips25_sap3/net262 ),
    .A2(\heichips25_sap3/net230 ));
 sg13g2_a221oi_1 \heichips25_sap3/_2278_  (.B2(\heichips25_sap3/net262 ),
    .C1(\heichips25_sap3/_1574_ ),
    .B1(\heichips25_sap3/_1662_ ),
    .A1(\heichips25_sap3/_1537_ ),
    .Y(\heichips25_sap3/_1699_ ),
    .A2(\heichips25_sap3/_1555_ ));
 sg13g2_and4_1 \heichips25_sap3/_2279_  (.A(\heichips25_sap3/_1659_ ),
    .B(\heichips25_sap3/_1660_ ),
    .C(\heichips25_sap3/_1698_ ),
    .D(\heichips25_sap3/_1699_ ),
    .X(\heichips25_sap3/_1700_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2280_  (.Y(\heichips25_sap3/_1701_ ),
    .B1(\heichips25_sap3/_1700_ ),
    .B2(\heichips25_sap3/_1564_ ),
    .A2(\heichips25_sap3/_1696_ ),
    .A1(\heichips25_sap3/_1539_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2281_  (.Y(\heichips25_sap3/_1702_ ),
    .A(\heichips25_sap3/net270 ),
    .B(\heichips25_sap3/_1617_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2282_  (.Y(\heichips25_sap3/_1703_ ),
    .A(\heichips25_sap3/_1629_ ),
    .B(\heichips25_sap3/_1702_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2283_  (.A(\heichips25_sap3/_1364_ ),
    .B(\heichips25_sap3/_1621_ ),
    .C(\heichips25_sap3/_1645_ ),
    .Y(\heichips25_sap3/_1704_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2284_  (.A(\heichips25_sap3/_1701_ ),
    .B(\heichips25_sap3/_1703_ ),
    .C(\heichips25_sap3/_1704_ ),
    .Y(\heichips25_sap3/_1705_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2285_  (.B1(\heichips25_sap3/net223 ),
    .Y(\heichips25_sap3/_1706_ ),
    .A1(\heichips25_sap3/_1701_ ),
    .A2(\heichips25_sap3/_1703_ ));
 sg13g2_nand3b_1 \heichips25_sap3/_2286_  (.B(\heichips25_sap3/_1706_ ),
    .C(\heichips25_sap3/_1641_ ),
    .Y(\heichips25_sap3/_1707_ ),
    .A_N(\heichips25_sap3/_1705_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2287_  (.A1(\heichips25_sap3/net270 ),
    .A2(\heichips25_sap3/_1649_ ),
    .Y(\heichips25_sap3/_1708_ ),
    .B1(\heichips25_sap3/_1453_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2288_  (.Y(\heichips25_sap3/_1709_ ),
    .A(\heichips25_sap3/net270 ),
    .B(\heichips25_sap3/_1651_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2289_  (.Y(\heichips25_sap3/_1710_ ),
    .A(\heichips25_sap3/_1453_ ),
    .B(\heichips25_sap3/_1709_ ));
 sg13g2_nand3_1 \heichips25_sap3/_2290_  (.B(\heichips25_sap3/_1679_ ),
    .C(\heichips25_sap3/_1710_ ),
    .A(\heichips25_sap3/net241 ),
    .Y(\heichips25_sap3/_1711_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2291_  (.A1(\heichips25_sap3/_1707_ ),
    .A2(\heichips25_sap3/_1708_ ),
    .Y(\heichips25_sap3/_1712_ ),
    .B1(\heichips25_sap3/_1711_ ));
 sg13g2_a21o_1 \heichips25_sap3/_2292_  (.A2(\heichips25_sap3/_1708_ ),
    .A1(\heichips25_sap3/_1707_ ),
    .B1(\heichips25_sap3/_1711_ ),
    .X(\heichips25_sap3/_1713_ ));
 sg13g2_nand3_1 \heichips25_sap3/_2293_  (.B(\heichips25_sap3/net227 ),
    .C(\heichips25_sap3/_1613_ ),
    .A(\heichips25_sap3/net273 ),
    .Y(\heichips25_sap3/_1714_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2294_  (.Y(\heichips25_sap3/_1715_ ),
    .A(\heichips25_sap3/net248 ),
    .B(\heichips25_sap3/_1714_ ));
 sg13g2_nand4_1 \heichips25_sap3/_2295_  (.B(\heichips25_sap3/_1491_ ),
    .C(\heichips25_sap3/_1538_ ),
    .A(\heichips25_sap3/net256 ),
    .Y(\heichips25_sap3/_1716_ ),
    .D(\heichips25_sap3/_1568_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2296_  (.A(\heichips25_sap3/_1435_ ),
    .B(\heichips25_sap3/_1613_ ),
    .Y(\heichips25_sap3/_1717_ ));
 sg13g2_nor4_1 \heichips25_sap3/_2297_  (.A(\heichips25_sap3/_1476_ ),
    .B(\heichips25_sap3/_1614_ ),
    .C(\heichips25_sap3/_1623_ ),
    .D(\heichips25_sap3/_1717_ ),
    .Y(\heichips25_sap3/_1718_ ));
 sg13g2_or4_1 \heichips25_sap3/_2298_  (.A(\heichips25_sap3/_1476_ ),
    .B(\heichips25_sap3/_1614_ ),
    .C(\heichips25_sap3/_1623_ ),
    .D(\heichips25_sap3/_1717_ ),
    .X(\heichips25_sap3/_1719_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2299_  (.A1(\heichips25_sap3/_1450_ ),
    .A2(\heichips25_sap3/_1718_ ),
    .Y(\heichips25_sap3/_1720_ ),
    .B1(\heichips25_sap3/_1616_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2300_  (.A(\heichips25_sap3/_1363_ ),
    .B(\heichips25_sap3/_1441_ ),
    .Y(\heichips25_sap3/_1721_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2301_  (.Y(\heichips25_sap3/_1722_ ),
    .A(\heichips25_sap3/net264 ),
    .B(\heichips25_sap3/net256 ));
 sg13g2_nor2_1 \heichips25_sap3/_2302_  (.A(\heichips25_sap3/net234 ),
    .B(\heichips25_sap3/_1722_ ),
    .Y(\heichips25_sap3/_1723_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2303_  (.A(\heichips25_sap3/_1536_ ),
    .B(\heichips25_sap3/_1572_ ),
    .Y(\heichips25_sap3/_1724_ ));
 sg13g2_nand3_1 \heichips25_sap3/_2304_  (.B(\heichips25_sap3/net245 ),
    .C(\heichips25_sap3/_1551_ ),
    .A(\heichips25_sap3/_1463_ ),
    .Y(\heichips25_sap3/_1725_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2305_  (.A(\heichips25_sap3/net264 ),
    .B(\heichips25_sap3/_1725_ ),
    .Y(\heichips25_sap3/_1726_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2306_  (.A(\heichips25_sap3/_1462_ ),
    .B(\heichips25_sap3/_1518_ ),
    .Y(\heichips25_sap3/_1727_ ));
 sg13g2_nor4_1 \heichips25_sap3/_2307_  (.A(\heichips25_sap3/_1599_ ),
    .B(\heichips25_sap3/net218 ),
    .C(\heichips25_sap3/_1726_ ),
    .D(\heichips25_sap3/_1727_ ),
    .Y(\heichips25_sap3/_1728_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2308_  (.Y(\heichips25_sap3/_1729_ ),
    .B1(\heichips25_sap3/_1723_ ),
    .B2(\heichips25_sap3/_1618_ ),
    .A2(\heichips25_sap3/_1720_ ),
    .A1(\heichips25_sap3/net272 ));
 sg13g2_nand4_1 \heichips25_sap3/_2309_  (.B(\heichips25_sap3/_1716_ ),
    .C(\heichips25_sap3/_1728_ ),
    .A(\heichips25_sap3/_1454_ ),
    .Y(\heichips25_sap3/_1730_ ),
    .D(\heichips25_sap3/_1729_ ));
 sg13g2_and2_1 \heichips25_sap3/_2310_  (.A(\heichips25_sap3/_1715_ ),
    .B(\heichips25_sap3/_1730_ ),
    .X(\heichips25_sap3/_1731_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2311_  (.Y(\heichips25_sap3/_1732_ ),
    .A(\heichips25_sap3/_1715_ ),
    .B(\heichips25_sap3/_1730_ ));
 sg13g2_nor4_1 \heichips25_sap3/_2312_  (.A(\heichips25_sap3/_1680_ ),
    .B(\heichips25_sap3/_1693_ ),
    .C(\heichips25_sap3/_1712_ ),
    .D(\heichips25_sap3/_1731_ ),
    .Y(\heichips25_sap3/_1733_ ));
 sg13g2_nand3_1 \heichips25_sap3/_2313_  (.B(\heichips25_sap3/_1713_ ),
    .C(\heichips25_sap3/_1732_ ),
    .A(\heichips25_sap3/_1695_ ),
    .Y(\heichips25_sap3/_1734_ ));
 sg13g2_nor4_1 \heichips25_sap3/_2314_  (.A(\heichips25_sap3/_1680_ ),
    .B(\heichips25_sap3/_1693_ ),
    .C(\heichips25_sap3/_1712_ ),
    .D(\heichips25_sap3/_1732_ ),
    .Y(\heichips25_sap3/_1735_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_2315_  (.B2(\heichips25_sap3/_1730_ ),
    .C1(\heichips25_sap3/_1711_ ),
    .B1(\heichips25_sap3/_1715_ ),
    .A1(\heichips25_sap3/_1708_ ),
    .Y(\heichips25_sap3/_1736_ ),
    .A2(\heichips25_sap3/_1707_ ));
 sg13g2_and2_1 \heichips25_sap3/_2316_  (.A(\heichips25_sap3/_1695_ ),
    .B(\heichips25_sap3/_1736_ ),
    .X(\heichips25_sap3/_1737_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2317_  (.Y(\heichips25_sap3/_1738_ ),
    .B1(\heichips25_sap3/net85 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][7] ),
    .A2(\heichips25_sap3/net87 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][7] ));
 sg13g2_nor4_1 \heichips25_sap3/_2318_  (.A(\heichips25_sap3/_1680_ ),
    .B(\heichips25_sap3/_1693_ ),
    .C(\heichips25_sap3/_1713_ ),
    .D(\heichips25_sap3/_1732_ ),
    .Y(\heichips25_sap3/_1739_ ));
 sg13g2_and3_1 \heichips25_sap3/_2319_  (.X(\heichips25_sap3/_1740_ ),
    .A(\heichips25_sap3/_1680_ ),
    .B(\heichips25_sap3/_1713_ ),
    .C(\heichips25_sap3/_1732_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2320_  (.A(\heichips25_sap3/_1694_ ),
    .B(\heichips25_sap3/_1713_ ),
    .C(\heichips25_sap3/_1732_ ),
    .Y(\heichips25_sap3/_1741_ ));
 sg13g2_nand3_1 \heichips25_sap3/_2321_  (.B(\heichips25_sap3/_1712_ ),
    .C(\heichips25_sap3/_1731_ ),
    .A(\heichips25_sap3/_1693_ ),
    .Y(\heichips25_sap3/_1742_ ));
 sg13g2_and2_1 \heichips25_sap3/_2322_  (.A(\heichips25_sap3/_1693_ ),
    .B(\heichips25_sap3/_1736_ ),
    .X(\heichips25_sap3/_1743_ ));
 sg13g2_and2_1 \heichips25_sap3/_2323_  (.A(\heichips25_sap3/_1680_ ),
    .B(\heichips25_sap3/_1736_ ),
    .X(\heichips25_sap3/_1744_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2324_  (.A(\heichips25_sap3/_1694_ ),
    .B(\heichips25_sap3/_1712_ ),
    .C(\heichips25_sap3/_1731_ ),
    .Y(\heichips25_sap3/_1745_ ));
 sg13g2_and3_1 \heichips25_sap3/_2325_  (.X(\heichips25_sap3/_1746_ ),
    .A(\heichips25_sap3/_1680_ ),
    .B(\heichips25_sap3/_1713_ ),
    .C(\heichips25_sap3/_1731_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_2326_  (.B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][7] ),
    .C1(\heichips25_sap3/net90 ),
    .B1(\heichips25_sap3/net75 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][7] ),
    .Y(\heichips25_sap3/_1747_ ),
    .A2(\heichips25_sap3/net77 ));
 sg13g2_a22oi_1 \heichips25_sap3/_2327_  (.Y(\heichips25_sap3/_1748_ ),
    .B1(\heichips25_sap3/net73 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][7] ),
    .A2(\heichips25_sap3/net83 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][7] ));
 sg13g2_a22oi_1 \heichips25_sap3/_2328_  (.Y(\heichips25_sap3/_1749_ ),
    .B1(\heichips25_sap3/net79 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][7] ),
    .A2(\heichips25_sap3/net81 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][7] ));
 sg13g2_a22oi_1 \heichips25_sap3/_2329_  (.Y(\heichips25_sap3/_1750_ ),
    .B1(\heichips25_sap3/net71 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][7] ),
    .A2(\heichips25_sap3/net216 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][7] ));
 sg13g2_and4_1 \heichips25_sap3/_2330_  (.A(\heichips25_sap3/_1738_ ),
    .B(\heichips25_sap3/_1748_ ),
    .C(\heichips25_sap3/_1749_ ),
    .D(\heichips25_sap3/_1750_ ),
    .X(\heichips25_sap3/_1751_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_2331_  (.B2(\heichips25_sap3/_1751_ ),
    .C1(\heichips25_sap3/_1654_ ),
    .B1(\heichips25_sap3/_1747_ ),
    .A1(\heichips25_sap3/_1420_ ),
    .Y(\heichips25_sap3/_1752_ ),
    .A2(\heichips25_sap3/net90 ));
 sg13g2_a21oi_1 \heichips25_sap3/_2332_  (.A1(\heichips25_sap3/net249 ),
    .A2(\heichips25_sap3/net225 ),
    .Y(\heichips25_sap3/_1753_ ),
    .B1(\heichips25_sap3/_1455_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2333_  (.A(\heichips25_sap3/net244 ),
    .B(\heichips25_sap3/_1530_ ),
    .C(\heichips25_sap3/_1531_ ),
    .Y(\heichips25_sap3/_1754_ ));
 sg13g2_nand3_1 \heichips25_sap3/_2334_  (.B(\heichips25_sap3/net242 ),
    .C(\heichips25_sap3/_1549_ ),
    .A(\heichips25_sap3/net266 ),
    .Y(\heichips25_sap3/_1755_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2335_  (.Y(\heichips25_sap3/_1756_ ),
    .B1(\heichips25_sap3/_1755_ ),
    .B2(\heichips25_sap3/_1486_ ),
    .A2(\heichips25_sap3/_1754_ ),
    .A1(\heichips25_sap3/_1685_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2336_  (.B1(\heichips25_sap3/_1486_ ),
    .Y(\heichips25_sap3/_1757_ ),
    .A1(\heichips25_sap3/_1363_ ),
    .A2(\heichips25_sap3/_1553_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2337_  (.Y(\heichips25_sap3/_1758_ ),
    .A(\heichips25_sap3/net245 ),
    .B(\heichips25_sap3/_1757_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2338_  (.A(\heichips25_sap3/_1486_ ),
    .B(\heichips25_sap3/_1495_ ),
    .Y(\heichips25_sap3/_1759_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2339_  (.A1(\heichips25_sap3/net227 ),
    .A2(\heichips25_sap3/_1623_ ),
    .Y(\heichips25_sap3/_1760_ ),
    .B1(\heichips25_sap3/net223 ));
 sg13g2_nand3_1 \heichips25_sap3/_2340_  (.B(\heichips25_sap3/_1515_ ),
    .C(\heichips25_sap3/_1605_ ),
    .A(\heichips25_sap3/net264 ),
    .Y(\heichips25_sap3/_1761_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2341_  (.A(\heichips25_sap3/_1475_ ),
    .B(\heichips25_sap3/net225 ),
    .Y(\heichips25_sap3/_1762_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2342_  (.A(\heichips25_sap3/_1759_ ),
    .B(\heichips25_sap3/_1762_ ),
    .Y(\heichips25_sap3/_1763_ ));
 sg13g2_nand4_1 \heichips25_sap3/_2343_  (.B(\heichips25_sap3/_1760_ ),
    .C(\heichips25_sap3/_1761_ ),
    .A(\heichips25_sap3/_1758_ ),
    .Y(\heichips25_sap3/_1764_ ),
    .D(\heichips25_sap3/_1763_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2344_  (.A1(\heichips25_sap3/net224 ),
    .A2(\heichips25_sap3/_1709_ ),
    .Y(\heichips25_sap3/_1765_ ),
    .B1(\heichips25_sap3/net220 ));
 sg13g2_o21ai_1 \heichips25_sap3/_2345_  (.B1(\heichips25_sap3/_1765_ ),
    .Y(\heichips25_sap3/_1766_ ),
    .A1(\heichips25_sap3/_1756_ ),
    .A2(\heichips25_sap3/_1764_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2346_  (.Y(\heichips25_sap3/_1767_ ),
    .A(\heichips25_sap3/_1472_ ),
    .B(\heichips25_sap3/net227 ));
 sg13g2_nand3_1 \heichips25_sap3/_2347_  (.B(\heichips25_sap3/_1766_ ),
    .C(\heichips25_sap3/_1767_ ),
    .A(\heichips25_sap3/_1452_ ),
    .Y(\heichips25_sap3/_1768_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2348_  (.Y(\heichips25_sap3/_1769_ ),
    .A(\heichips25_sap3/_1753_ ),
    .B(\heichips25_sap3/_1768_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2349_  (.Y(\heichips25_sap3/_1770_ ),
    .A(\heichips25_sap3/net231 ),
    .B(\heichips25_sap3/_1769_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2350_  (.Y(\heichips25_sap3/_1771_ ),
    .A(net10),
    .B(\heichips25_sap3/_1770_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2351_  (.A(\heichips25_sap3/_1454_ ),
    .B(\heichips25_sap3/net226 ),
    .C(\heichips25_sap3/_1613_ ),
    .Y(\heichips25_sap3/_1772_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2352_  (.A(\heichips25_sap3/_1480_ ),
    .B(\heichips25_sap3/_1619_ ),
    .Y(\heichips25_sap3/_1773_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2353_  (.Y(\heichips25_sap3/_1774_ ),
    .B1(\heichips25_sap3/_1605_ ),
    .B2(\heichips25_sap3/_1515_ ),
    .A2(\heichips25_sap3/_1549_ ),
    .A1(\heichips25_sap3/net242 ));
 sg13g2_or2_1 \heichips25_sap3/_2354_  (.X(\heichips25_sap3/_1775_ ),
    .B(\heichips25_sap3/_1774_ ),
    .A(\heichips25_sap3/net266 ));
 sg13g2_a21oi_1 \heichips25_sap3/_2355_  (.A1(\heichips25_sap3/_1517_ ),
    .A2(\heichips25_sap3/_1549_ ),
    .Y(\heichips25_sap3/_1776_ ),
    .B1(\heichips25_sap3/net223 ));
 sg13g2_nor3_1 \heichips25_sap3/_2356_  (.A(\heichips25_sap3/net256 ),
    .B(\heichips25_sap3/_1480_ ),
    .C(\heichips25_sap3/_1492_ ),
    .Y(\heichips25_sap3/_1777_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2357_  (.A1(\heichips25_sap3/net229 ),
    .A2(\heichips25_sap3/_1550_ ),
    .Y(\heichips25_sap3/_1778_ ),
    .B1(\heichips25_sap3/_1518_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2358_  (.A(\heichips25_sap3/net223 ),
    .B(\heichips25_sap3/_1777_ ),
    .C(\heichips25_sap3/_1778_ ),
    .Y(\heichips25_sap3/_1779_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2359_  (.Y(\heichips25_sap3/_1780_ ),
    .A(\heichips25_sap3/_1775_ ),
    .B(\heichips25_sap3/_1779_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2360_  (.B1(\heichips25_sap3/_1780_ ),
    .Y(\heichips25_sap3/_1781_ ),
    .A1(\heichips25_sap3/_1621_ ),
    .A2(\heichips25_sap3/_1773_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2361_  (.A(\heichips25_sap3/_1458_ ),
    .B(\heichips25_sap3/_1460_ ),
    .C(\heichips25_sap3/_1613_ ),
    .Y(\heichips25_sap3/_1782_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2362_  (.Y(\heichips25_sap3/_1783_ ),
    .A(\heichips25_sap3/_1472_ ),
    .B(\heichips25_sap3/_1496_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2363_  (.Y(\heichips25_sap3/_1784_ ),
    .A(\heichips25_sap3/net220 ),
    .B(\heichips25_sap3/_1783_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2364_  (.A1(\heichips25_sap3/_1449_ ),
    .A2(\heichips25_sap3/_1782_ ),
    .Y(\heichips25_sap3/_1785_ ),
    .B1(\heichips25_sap3/_1784_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2365_  (.A1(\heichips25_sap3/_1641_ ),
    .A2(\heichips25_sap3/_1781_ ),
    .Y(\heichips25_sap3/_1786_ ),
    .B1(\heichips25_sap3/_1785_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2366_  (.A1(\heichips25_sap3/_1454_ ),
    .A2(\heichips25_sap3/_1786_ ),
    .Y(\heichips25_sap3/_1787_ ),
    .B1(\heichips25_sap3/_1772_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2367_  (.A(\heichips25_sap3/net256 ),
    .B(\heichips25_sap3/_1492_ ),
    .C(\heichips25_sap3/_1569_ ),
    .Y(\heichips25_sap3/_1788_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2368_  (.Y(\heichips25_sap3/_1789_ ),
    .A(\heichips25_sap3/sap_3_inst.alu_flags[7] ),
    .B(\heichips25_sap3/_1788_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2369_  (.Y(\heichips25_sap3/_1790_ ),
    .A(\heichips25_sap3/net155 ),
    .B(\heichips25_sap3/_1789_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2370_  (.B1(\heichips25_sap3/_1790_ ),
    .Y(\heichips25_sap3/_1791_ ),
    .A1(\heichips25_sap3/net274 ),
    .A2(\heichips25_sap3/net155 ));
 sg13g2_nand2_1 \heichips25_sap3/_2371_  (.Y(\heichips25_sap3/_1792_ ),
    .A(\heichips25_sap3/_1771_ ),
    .B(\heichips25_sap3/_1791_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2372_  (.Y(\heichips25_sap3/_1793_ ),
    .B1(\heichips25_sap3/net72 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][7] ),
    .A2(\heichips25_sap3/net85 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][7] ));
 sg13g2_a22oi_1 \heichips25_sap3/_2373_  (.Y(\heichips25_sap3/_1794_ ),
    .B1(\heichips25_sap3/net75 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][7] ),
    .A2(\heichips25_sap3/net81 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][7] ));
 sg13g2_and2_1 \heichips25_sap3/_2374_  (.A(\heichips25_sap3/_1793_ ),
    .B(\heichips25_sap3/_1794_ ),
    .X(\heichips25_sap3/_1795_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_2375_  (.B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][7] ),
    .C1(\heichips25_sap3/net79 ),
    .B1(\heichips25_sap3/net84 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][7] ),
    .Y(\heichips25_sap3/_1796_ ),
    .A2(\heichips25_sap3/net216 ));
 sg13g2_a22oi_1 \heichips25_sap3/_2376_  (.Y(\heichips25_sap3/_1797_ ),
    .B1(\heichips25_sap3/net73 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][7] ),
    .A2(\heichips25_sap3/net90 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][7] ));
 sg13g2_a22oi_1 \heichips25_sap3/_2377_  (.Y(\heichips25_sap3/_1798_ ),
    .B1(\heichips25_sap3/net77 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][7] ),
    .A2(\heichips25_sap3/net87 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][7] ));
 sg13g2_and3_1 \heichips25_sap3/_2378_  (.X(\heichips25_sap3/_1799_ ),
    .A(\heichips25_sap3/_1796_ ),
    .B(\heichips25_sap3/_1797_ ),
    .C(\heichips25_sap3/_1798_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2379_  (.A1(\heichips25_sap3/_1795_ ),
    .A2(\heichips25_sap3/_1799_ ),
    .Y(\heichips25_sap3/_1800_ ),
    .B1(\heichips25_sap3/net66 ));
 sg13g2_or3_1 \heichips25_sap3/_2380_  (.A(\heichips25_sap3/_1752_ ),
    .B(\heichips25_sap3/_1792_ ),
    .C(\heichips25_sap3/_1800_ ),
    .X(\uio_out_sap3[7] ));
 sg13g2_nor3_1 \heichips25_sap3/_2381_  (.A(\heichips25_sap3/_1442_ ),
    .B(\heichips25_sap3/_1495_ ),
    .C(\heichips25_sap3/net226 ),
    .Y(\heichips25_sap3/_1801_ ));
 sg13g2_nand3_1 \heichips25_sap3/_2382_  (.B(\heichips25_sap3/_1494_ ),
    .C(\heichips25_sap3/net227 ),
    .A(\heichips25_sap3/_1441_ ),
    .Y(\heichips25_sap3/_1802_ ));
 sg13g2_mux2_1 \heichips25_sap3/_2383_  (.A0(\heichips25_sap3/sap_3_inst.alu_flags[7] ),
    .A1(net47),
    .S(\heichips25_sap3/net215 ),
    .X(\heichips25_sap3/_0038_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2384_  (.A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[0][6] ),
    .B(\heichips25_sap3/_1734_ ),
    .Y(\heichips25_sap3/_1803_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2385_  (.Y(\heichips25_sap3/_1804_ ),
    .B1(\heichips25_sap3/net73 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][6] ),
    .A2(\heichips25_sap3/net77 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][6] ));
 sg13g2_a22oi_1 \heichips25_sap3/_2386_  (.Y(\heichips25_sap3/_1805_ ),
    .B1(\heichips25_sap3/net72 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][6] ),
    .A2(\heichips25_sap3/net216 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][6] ));
 sg13g2_a22oi_1 \heichips25_sap3/_2387_  (.Y(\heichips25_sap3/_1806_ ),
    .B1(\heichips25_sap3/net81 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][6] ),
    .A2(\heichips25_sap3/net87 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][6] ));
 sg13g2_a22oi_1 \heichips25_sap3/_2388_  (.Y(\heichips25_sap3/_1807_ ),
    .B1(\heichips25_sap3/net80 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][6] ),
    .A2(\heichips25_sap3/net84 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][6] ));
 sg13g2_nand2_1 \heichips25_sap3/_2389_  (.Y(\heichips25_sap3/_1808_ ),
    .A(\heichips25_sap3/_1806_ ),
    .B(\heichips25_sap3/_1807_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2390_  (.Y(\heichips25_sap3/_1809_ ),
    .B1(\heichips25_sap3/net75 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][6] ),
    .A2(\heichips25_sap3/net85 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][6] ));
 sg13g2_nand4_1 \heichips25_sap3/_2391_  (.B(\heichips25_sap3/_1804_ ),
    .C(\heichips25_sap3/_1805_ ),
    .A(\heichips25_sap3/_1734_ ),
    .Y(\heichips25_sap3/_1810_ ),
    .D(\heichips25_sap3/_1809_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2392_  (.A(\heichips25_sap3/_1808_ ),
    .B(\heichips25_sap3/_1810_ ),
    .Y(\heichips25_sap3/_1811_ ));
 sg13g2_or3_1 \heichips25_sap3/_2393_  (.A(\heichips25_sap3/_1654_ ),
    .B(\heichips25_sap3/_1803_ ),
    .C(\heichips25_sap3/_1811_ ),
    .X(\heichips25_sap3/_1812_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2394_  (.Y(\heichips25_sap3/_1813_ ),
    .A(net9),
    .B(\heichips25_sap3/_1770_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2395_  (.Y(\heichips25_sap3/_1814_ ),
    .A(\heichips25_sap3/sap_3_inst.alu_flags[6] ),
    .B(\heichips25_sap3/_1788_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2396_  (.Y(\heichips25_sap3/_1815_ ),
    .A(\heichips25_sap3/net155 ),
    .B(\heichips25_sap3/_1814_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2397_  (.B1(\heichips25_sap3/_1815_ ),
    .Y(\heichips25_sap3/_1816_ ),
    .A1(\heichips25_sap3/net277 ),
    .A2(\heichips25_sap3/net155 ));
 sg13g2_a22oi_1 \heichips25_sap3/_2398_  (.Y(\heichips25_sap3/_1817_ ),
    .B1(\heichips25_sap3/net75 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][6] ),
    .A2(\heichips25_sap3/net84 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][6] ));
 sg13g2_a22oi_1 \heichips25_sap3/_2399_  (.Y(\heichips25_sap3/_1818_ ),
    .B1(\heichips25_sap3/net77 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][6] ),
    .A2(\heichips25_sap3/net90 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][6] ));
 sg13g2_a22oi_1 \heichips25_sap3/_2400_  (.Y(\heichips25_sap3/_1819_ ),
    .B1(\heichips25_sap3/net73 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][6] ),
    .A2(\heichips25_sap3/net81 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][6] ));
 sg13g2_a22oi_1 \heichips25_sap3/_2401_  (.Y(\heichips25_sap3/_1820_ ),
    .B1(\heichips25_sap3/net72 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][6] ),
    .A2(\heichips25_sap3/net216 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][6] ));
 sg13g2_nand4_1 \heichips25_sap3/_2402_  (.B(\heichips25_sap3/_1817_ ),
    .C(\heichips25_sap3/_1819_ ),
    .A(\heichips25_sap3/_1742_ ),
    .Y(\heichips25_sap3/_1821_ ),
    .D(\heichips25_sap3/_1820_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_2403_  (.B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][6] ),
    .C1(\heichips25_sap3/_1821_ ),
    .B1(\heichips25_sap3/net85 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][6] ),
    .Y(\heichips25_sap3/_1822_ ),
    .A2(\heichips25_sap3/net87 ));
 sg13g2_a21o_1 \heichips25_sap3/_2404_  (.A2(\heichips25_sap3/_1822_ ),
    .A1(\heichips25_sap3/_1818_ ),
    .B1(\heichips25_sap3/net66 ),
    .X(\heichips25_sap3/_1823_ ));
 sg13g2_nand4_1 \heichips25_sap3/_2405_  (.B(\heichips25_sap3/_1813_ ),
    .C(\heichips25_sap3/_1816_ ),
    .A(\heichips25_sap3/_1823_ ),
    .Y(\uio_out_sap3[6] ),
    .D(\heichips25_sap3/_1812_ ));
 sg13g2_mux2_1 \heichips25_sap3/_2406_  (.A0(\heichips25_sap3/sap_3_inst.alu_flags[6] ),
    .A1(net43),
    .S(\heichips25_sap3/net215 ),
    .X(\heichips25_sap3/_0037_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2407_  (.Y(\heichips25_sap3/_1824_ ),
    .B1(\heichips25_sap3/net80 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][5] ),
    .A2(\heichips25_sap3/net86 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][5] ));
 sg13g2_a22oi_1 \heichips25_sap3/_2408_  (.Y(\heichips25_sap3/_1825_ ),
    .B1(\heichips25_sap3/net84 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][5] ),
    .A2(\heichips25_sap3/net87 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][5] ));
 sg13g2_a22oi_1 \heichips25_sap3/_2409_  (.Y(\heichips25_sap3/_1826_ ),
    .B1(\heichips25_sap3/net75 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][5] ),
    .A2(\heichips25_sap3/net81 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][5] ));
 sg13g2_and2_1 \heichips25_sap3/_2410_  (.A(\heichips25_sap3/_1825_ ),
    .B(\heichips25_sap3/_1826_ ),
    .X(\heichips25_sap3/_1827_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2411_  (.Y(\heichips25_sap3/_1828_ ),
    .B1(\heichips25_sap3/net72 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][5] ),
    .A2(\heichips25_sap3/net217 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][5] ));
 sg13g2_a22oi_1 \heichips25_sap3/_2412_  (.Y(\heichips25_sap3/_1829_ ),
    .B1(\heichips25_sap3/_1745_ ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][5] ),
    .A2(\heichips25_sap3/_1743_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][5] ));
 sg13g2_and4_1 \heichips25_sap3/_2413_  (.A(\heichips25_sap3/_1734_ ),
    .B(\heichips25_sap3/_1824_ ),
    .C(\heichips25_sap3/_1828_ ),
    .D(\heichips25_sap3/_1829_ ),
    .X(\heichips25_sap3/_1830_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_2414_  (.B2(\heichips25_sap3/_1830_ ),
    .C1(\heichips25_sap3/_1654_ ),
    .B1(\heichips25_sap3/_1827_ ),
    .A1(\heichips25_sap3/_1404_ ),
    .Y(\heichips25_sap3/_1831_ ),
    .A2(\heichips25_sap3/net91 ));
 sg13g2_nand2_1 \heichips25_sap3/_2415_  (.Y(\heichips25_sap3/_1832_ ),
    .A(\heichips25_sap3/sap_3_inst.alu_flags[5] ),
    .B(\heichips25_sap3/_1788_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2416_  (.Y(\heichips25_sap3/_1833_ ),
    .A(\heichips25_sap3/net155 ),
    .B(\heichips25_sap3/_1832_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2417_  (.B1(\heichips25_sap3/_1833_ ),
    .Y(\heichips25_sap3/_1834_ ),
    .A1(\heichips25_sap3/net279 ),
    .A2(\heichips25_sap3/net155 ));
 sg13g2_nand2_1 \heichips25_sap3/_2418_  (.Y(\heichips25_sap3/_1835_ ),
    .A(net8),
    .B(\heichips25_sap3/_1770_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2419_  (.Y(\heichips25_sap3/_1836_ ),
    .A(\heichips25_sap3/_1834_ ),
    .B(\heichips25_sap3/_1835_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2420_  (.Y(\heichips25_sap3/_1837_ ),
    .B1(\heichips25_sap3/net78 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][5] ),
    .A2(\heichips25_sap3/net86 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][5] ));
 sg13g2_a22oi_1 \heichips25_sap3/_2421_  (.Y(\heichips25_sap3/_1838_ ),
    .B1(\heichips25_sap3/net72 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][5] ),
    .A2(\heichips25_sap3/_1744_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][5] ));
 sg13g2_and2_1 \heichips25_sap3/_2422_  (.A(\heichips25_sap3/_1837_ ),
    .B(\heichips25_sap3/_1838_ ),
    .X(\heichips25_sap3/_1839_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_2423_  (.B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][5] ),
    .C1(\heichips25_sap3/net80 ),
    .B1(\heichips25_sap3/net74 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][5] ),
    .Y(\heichips25_sap3/_1840_ ),
    .A2(\heichips25_sap3/net217 ));
 sg13g2_a22oi_1 \heichips25_sap3/_2424_  (.Y(\heichips25_sap3/_1841_ ),
    .B1(\heichips25_sap3/_1740_ ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][5] ),
    .A2(\heichips25_sap3/net88 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][5] ));
 sg13g2_a22oi_1 \heichips25_sap3/_2425_  (.Y(\heichips25_sap3/_1842_ ),
    .B1(\heichips25_sap3/net84 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][5] ),
    .A2(\heichips25_sap3/net91 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][5] ));
 sg13g2_and3_1 \heichips25_sap3/_2426_  (.X(\heichips25_sap3/_1843_ ),
    .A(\heichips25_sap3/_1840_ ),
    .B(\heichips25_sap3/_1841_ ),
    .C(\heichips25_sap3/_1842_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2427_  (.A1(\heichips25_sap3/_1839_ ),
    .A2(\heichips25_sap3/_1843_ ),
    .Y(\heichips25_sap3/_1844_ ),
    .B1(\heichips25_sap3/net66 ));
 sg13g2_or3_1 \heichips25_sap3/_2428_  (.A(\heichips25_sap3/_1831_ ),
    .B(\heichips25_sap3/_1836_ ),
    .C(\heichips25_sap3/_1844_ ),
    .X(\uio_out_sap3[5] ));
 sg13g2_mux2_1 \heichips25_sap3/_2429_  (.A0(\heichips25_sap3/sap_3_inst.alu_flags[5] ),
    .A1(\uio_out_sap3[5] ),
    .S(\heichips25_sap3/net215 ),
    .X(\heichips25_sap3/_0036_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2430_  (.Y(\heichips25_sap3/_1845_ ),
    .B1(\heichips25_sap3/net85 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][4] ),
    .A2(\heichips25_sap3/net87 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][4] ));
 sg13g2_a22oi_1 \heichips25_sap3/_2431_  (.Y(\heichips25_sap3/_1846_ ),
    .B1(\heichips25_sap3/net75 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][4] ),
    .A2(\heichips25_sap3/net81 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][4] ));
 sg13g2_a22oi_1 \heichips25_sap3/_2432_  (.Y(\heichips25_sap3/_1847_ ),
    .B1(\heichips25_sap3/net80 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][4] ),
    .A2(\heichips25_sap3/net84 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][4] ));
 sg13g2_and2_1 \heichips25_sap3/_2433_  (.A(\heichips25_sap3/_1845_ ),
    .B(\heichips25_sap3/_1847_ ),
    .X(\heichips25_sap3/_1848_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2434_  (.Y(\heichips25_sap3/_1849_ ),
    .B1(\heichips25_sap3/net72 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][4] ),
    .A2(\heichips25_sap3/net217 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][4] ));
 sg13g2_a22oi_1 \heichips25_sap3/_2435_  (.Y(\heichips25_sap3/_1850_ ),
    .B1(\heichips25_sap3/net73 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][4] ),
    .A2(\heichips25_sap3/net77 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][4] ));
 sg13g2_and4_1 \heichips25_sap3/_2436_  (.A(\heichips25_sap3/_1734_ ),
    .B(\heichips25_sap3/_1846_ ),
    .C(\heichips25_sap3/_1849_ ),
    .D(\heichips25_sap3/_1850_ ),
    .X(\heichips25_sap3/_1851_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_2437_  (.B2(\heichips25_sap3/_1851_ ),
    .C1(\heichips25_sap3/_1654_ ),
    .B1(\heichips25_sap3/_1848_ ),
    .A1(\heichips25_sap3/_1400_ ),
    .Y(\heichips25_sap3/_1852_ ),
    .A2(\heichips25_sap3/net90 ));
 sg13g2_or2_1 \heichips25_sap3/_2438_  (.X(\heichips25_sap3/_1853_ ),
    .B(\heichips25_sap3/net155 ),
    .A(\heichips25_sap3/net280 ));
 sg13g2_nand2_1 \heichips25_sap3/_2439_  (.Y(\heichips25_sap3/_1854_ ),
    .A(\heichips25_sap3/sap_3_inst.alu_flags[4] ),
    .B(\heichips25_sap3/_1788_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2440_  (.Y(\heichips25_sap3/_1855_ ),
    .A(\heichips25_sap3/net156 ),
    .B(\heichips25_sap3/_1854_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2441_  (.Y(\heichips25_sap3/_1856_ ),
    .B1(\heichips25_sap3/_1853_ ),
    .B2(\heichips25_sap3/_1855_ ),
    .A2(\heichips25_sap3/_1770_ ),
    .A1(net7));
 sg13g2_a22oi_1 \heichips25_sap3/_2442_  (.Y(\heichips25_sap3/_1857_ ),
    .B1(\heichips25_sap3/net75 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][4] ),
    .A2(\heichips25_sap3/net90 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][4] ));
 sg13g2_a22oi_1 \heichips25_sap3/_2443_  (.Y(\heichips25_sap3/_1858_ ),
    .B1(\heichips25_sap3/net73 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][4] ),
    .A2(\heichips25_sap3/net81 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][4] ));
 sg13g2_and2_1 \heichips25_sap3/_2444_  (.A(\heichips25_sap3/_1857_ ),
    .B(\heichips25_sap3/_1858_ ),
    .X(\heichips25_sap3/_1859_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_2445_  (.B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][4] ),
    .C1(\heichips25_sap3/net80 ),
    .B1(\heichips25_sap3/net72 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][4] ),
    .Y(\heichips25_sap3/_1860_ ),
    .A2(\heichips25_sap3/net217 ));
 sg13g2_a22oi_1 \heichips25_sap3/_2446_  (.Y(\heichips25_sap3/_1861_ ),
    .B1(\heichips25_sap3/net85 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][4] ),
    .A2(\heichips25_sap3/net87 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][4] ));
 sg13g2_a22oi_1 \heichips25_sap3/_2447_  (.Y(\heichips25_sap3/_1862_ ),
    .B1(\heichips25_sap3/net77 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][4] ),
    .A2(\heichips25_sap3/net84 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][4] ));
 sg13g2_and3_1 \heichips25_sap3/_2448_  (.X(\heichips25_sap3/_1863_ ),
    .A(\heichips25_sap3/_1860_ ),
    .B(\heichips25_sap3/_1861_ ),
    .C(\heichips25_sap3/_1862_ ));
 sg13g2_a21o_1 \heichips25_sap3/_2449_  (.A2(\heichips25_sap3/_1863_ ),
    .A1(\heichips25_sap3/_1859_ ),
    .B1(\heichips25_sap3/net66 ),
    .X(\heichips25_sap3/_1864_ ));
 sg13g2_nand3b_1 \heichips25_sap3/_2450_  (.B(\heichips25_sap3/_1856_ ),
    .C(\heichips25_sap3/_1864_ ),
    .Y(\uio_out_sap3[4] ),
    .A_N(\heichips25_sap3/_1852_ ));
 sg13g2_mux2_1 \heichips25_sap3/_2451_  (.A0(\heichips25_sap3/sap_3_inst.alu_flags[4] ),
    .A1(net46),
    .S(\heichips25_sap3/net215 ),
    .X(\heichips25_sap3/_0035_ ));
 sg13g2_nand3_1 \heichips25_sap3/_2452_  (.B(\heichips25_sap3/_1447_ ),
    .C(\heichips25_sap3/net230 ),
    .A(\heichips25_sap3/net259 ),
    .Y(\heichips25_sap3/_1865_ ));
 sg13g2_a21o_1 \heichips25_sap3/_2453_  (.A2(\heichips25_sap3/_1865_ ),
    .A1(\heichips25_sap3/net224 ),
    .B1(\heichips25_sap3/net221 ),
    .X(\heichips25_sap3/_1866_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2454_  (.A1(\heichips25_sap3/net238 ),
    .A2(\heichips25_sap3/_1643_ ),
    .Y(\heichips25_sap3/_1867_ ),
    .B1(\heichips25_sap3/net227 ));
 sg13g2_nor3_1 \heichips25_sap3/_2455_  (.A(\heichips25_sap3/_1619_ ),
    .B(\heichips25_sap3/net221 ),
    .C(\heichips25_sap3/_1867_ ),
    .Y(\heichips25_sap3/_1868_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2456_  (.A1(\heichips25_sap3/_1472_ ),
    .A2(\heichips25_sap3/net230 ),
    .Y(\heichips25_sap3/_1869_ ),
    .B1(\heichips25_sap3/_1868_ ));
 sg13g2_a21o_1 \heichips25_sap3/_2457_  (.A2(\heichips25_sap3/net230 ),
    .A1(\heichips25_sap3/_1472_ ),
    .B1(\heichips25_sap3/_1868_ ),
    .X(\heichips25_sap3/_1870_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2458_  (.A(\heichips25_sap3/net230 ),
    .B(\heichips25_sap3/_1559_ ),
    .Y(\heichips25_sap3/_1871_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2459_  (.A(\heichips25_sap3/_1518_ ),
    .B(\heichips25_sap3/_1871_ ),
    .Y(\heichips25_sap3/_1872_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2460_  (.A1(\heichips25_sap3/_1479_ ),
    .A2(\heichips25_sap3/_1623_ ),
    .Y(\heichips25_sap3/_1873_ ),
    .B1(\heichips25_sap3/_1872_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2461_  (.Y(\heichips25_sap3/_1874_ ),
    .B1(\heichips25_sap3/_1782_ ),
    .B2(\heichips25_sap3/_1361_ ),
    .A2(\heichips25_sap3/_1614_ ),
    .A1(\heichips25_sap3/net228 ));
 sg13g2_nand2_1 \heichips25_sap3/_2462_  (.Y(\heichips25_sap3/_1875_ ),
    .A(\heichips25_sap3/_1621_ ),
    .B(\heichips25_sap3/_1874_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2463_  (.A(\heichips25_sap3/net221 ),
    .B(\heichips25_sap3/_1875_ ),
    .Y(\heichips25_sap3/_1876_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2464_  (.Y(\heichips25_sap3/_1877_ ),
    .B1(\heichips25_sap3/_1873_ ),
    .B2(\heichips25_sap3/_1876_ ),
    .A2(\heichips25_sap3/_1869_ ),
    .A1(\heichips25_sap3/_1866_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2465_  (.A(\heichips25_sap3/net215 ),
    .B(\heichips25_sap3/_1877_ ),
    .Y(\heichips25_sap3/_1878_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2466_  (.B1(\heichips25_sap3/_1865_ ),
    .Y(\heichips25_sap3/_1879_ ),
    .A1(\heichips25_sap3/net224 ),
    .A2(\heichips25_sap3/_1874_ ));
 sg13g2_and2_1 \heichips25_sap3/_2467_  (.A(\heichips25_sap3/sap_3_inst.controller_inst.opcode[5] ),
    .B(\heichips25_sap3/_1879_ ),
    .X(\heichips25_sap3/_1880_ ));
 sg13g2_and2_1 \heichips25_sap3/_2468_  (.A(\heichips25_sap3/_1434_ ),
    .B(\heichips25_sap3/_1782_ ),
    .X(\heichips25_sap3/_1881_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2469_  (.Y(\heichips25_sap3/_1882_ ),
    .A(\heichips25_sap3/_1434_ ),
    .B(\heichips25_sap3/_1782_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2470_  (.Y(\heichips25_sap3/_1883_ ),
    .A(\heichips25_sap3/_1880_ ),
    .B(\heichips25_sap3/_1882_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2471_  (.Y(\heichips25_sap3/_1884_ ),
    .A(\heichips25_sap3/net263 ),
    .B(\heichips25_sap3/_1879_ ));
 sg13g2_nand3_1 \heichips25_sap3/_2472_  (.B(\heichips25_sap3/_1880_ ),
    .C(\heichips25_sap3/_1882_ ),
    .A(\heichips25_sap3/_1364_ ),
    .Y(\heichips25_sap3/_1885_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2473_  (.A(\heichips25_sap3/_1880_ ),
    .B(\heichips25_sap3/_1881_ ),
    .Y(\heichips25_sap3/_1886_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2474_  (.Y(\heichips25_sap3/_1887_ ),
    .A(\heichips25_sap3/_1869_ ),
    .B(\heichips25_sap3/_1886_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2475_  (.Y(\heichips25_sap3/_1888_ ),
    .A(\heichips25_sap3/sap_3_inst.controller_inst.opcode[4] ),
    .B(\heichips25_sap3/_1881_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2476_  (.A(\heichips25_sap3/_1619_ ),
    .B(\heichips25_sap3/_1714_ ),
    .Y(\heichips25_sap3/_1889_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2477_  (.A1(\heichips25_sap3/net265 ),
    .A2(\heichips25_sap3/_1879_ ),
    .Y(\heichips25_sap3/_1890_ ),
    .B1(\heichips25_sap3/net212 ));
 sg13g2_o21ai_1 \heichips25_sap3/_2478_  (.B1(\heichips25_sap3/_1890_ ),
    .Y(\heichips25_sap3/_1891_ ),
    .A1(\heichips25_sap3/_1518_ ),
    .A2(\heichips25_sap3/_1560_ ));
 sg13g2_nor2b_1 \heichips25_sap3/_2479_  (.A(\heichips25_sap3/_1884_ ),
    .B_N(\heichips25_sap3/net168 ),
    .Y(\heichips25_sap3/_1892_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_2480_  (.Y(\heichips25_sap3/_1893_ ),
    .B(\heichips25_sap3/net168 ),
    .A_N(\heichips25_sap3/_1884_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2481_  (.A(\heichips25_sap3/_1884_ ),
    .B(\heichips25_sap3/net168 ),
    .Y(\heichips25_sap3/_1894_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2482_  (.A(\heichips25_sap3/_1883_ ),
    .B(\heichips25_sap3/_1884_ ),
    .C(\heichips25_sap3/net168 ),
    .Y(\heichips25_sap3/_1895_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2483_  (.A(\heichips25_sap3/_1880_ ),
    .B(\heichips25_sap3/_1882_ ),
    .Y(\heichips25_sap3/_1896_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2484_  (.B1(\heichips25_sap3/_1893_ ),
    .Y(\heichips25_sap3/_1897_ ),
    .A1(\heichips25_sap3/net159 ),
    .A2(\heichips25_sap3/_1896_ ));
 sg13g2_and4_1 \heichips25_sap3/_2485_  (.A(\heichips25_sap3/_1885_ ),
    .B(\heichips25_sap3/_1887_ ),
    .C(\heichips25_sap3/_1888_ ),
    .D(\heichips25_sap3/_1897_ ),
    .X(\heichips25_sap3/_1898_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2486_  (.A(\heichips25_sap3/_1878_ ),
    .B(\heichips25_sap3/_1898_ ),
    .Y(\heichips25_sap3/_1899_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2487_  (.B1(\heichips25_sap3/net254 ),
    .Y(\heichips25_sap3/_1900_ ),
    .A1(\heichips25_sap3/_1878_ ),
    .A2(\heichips25_sap3/_1898_ ));
 sg13g2_and2_1 \heichips25_sap3/_2488_  (.A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][1] ),
    .B(\heichips25_sap3/net76 ),
    .X(\heichips25_sap3/_1901_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2489_  (.Y(\heichips25_sap3/_1902_ ),
    .B1(\heichips25_sap3/net74 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][1] ),
    .A2(\heichips25_sap3/net78 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][1] ));
 sg13g2_a22oi_1 \heichips25_sap3/_2490_  (.Y(\heichips25_sap3/_1903_ ),
    .B1(\heichips25_sap3/net86 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][1] ),
    .A2(\heichips25_sap3/net218 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][1] ));
 sg13g2_a221oi_1 \heichips25_sap3/_2491_  (.B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][1] ),
    .C1(\heichips25_sap3/_1901_ ),
    .B1(\heichips25_sap3/net71 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][1] ),
    .Y(\heichips25_sap3/_1904_ ),
    .A2(\heichips25_sap3/net79 ));
 sg13g2_a21oi_1 \heichips25_sap3/_2492_  (.A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][1] ),
    .A2(\heichips25_sap3/net88 ),
    .Y(\heichips25_sap3/_1905_ ),
    .B1(\heichips25_sap3/net89 ));
 sg13g2_a22oi_1 \heichips25_sap3/_2493_  (.Y(\heichips25_sap3/_1906_ ),
    .B1(\heichips25_sap3/net82 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][1] ),
    .A2(\heichips25_sap3/net83 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][1] ));
 sg13g2_and4_1 \heichips25_sap3/_2494_  (.A(\heichips25_sap3/_1902_ ),
    .B(\heichips25_sap3/_1903_ ),
    .C(\heichips25_sap3/_1905_ ),
    .D(\heichips25_sap3/_1906_ ),
    .X(\heichips25_sap3/_1907_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_2495_  (.B2(\heichips25_sap3/_1907_ ),
    .C1(\heichips25_sap3/_1654_ ),
    .B1(\heichips25_sap3/_1904_ ),
    .A1(\heichips25_sap3/_1385_ ),
    .Y(\heichips25_sap3/_1908_ ),
    .A2(\heichips25_sap3/net89 ));
 sg13g2_nand2_1 \heichips25_sap3/_2496_  (.Y(\heichips25_sap3/_1909_ ),
    .A(net4),
    .B(\heichips25_sap3/_1770_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2497_  (.Y(\heichips25_sap3/_1910_ ),
    .A(\heichips25_sap3/sap_3_inst.alu_flags[1] ),
    .B(\heichips25_sap3/_1788_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2498_  (.Y(\heichips25_sap3/_1911_ ),
    .A(\heichips25_sap3/net156 ),
    .B(\heichips25_sap3/_1910_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2499_  (.B1(\heichips25_sap3/_1911_ ),
    .Y(\heichips25_sap3/_1912_ ),
    .A1(\heichips25_sap3/net286 ),
    .A2(\heichips25_sap3/net156 ));
 sg13g2_nand2_1 \heichips25_sap3/_2500_  (.Y(\heichips25_sap3/_1913_ ),
    .A(\heichips25_sap3/_1909_ ),
    .B(\heichips25_sap3/_1912_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2501_  (.Y(\heichips25_sap3/_1914_ ),
    .B1(\heichips25_sap3/net71 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][1] ),
    .A2(\heichips25_sap3/net74 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][1] ));
 sg13g2_a22oi_1 \heichips25_sap3/_2502_  (.Y(\heichips25_sap3/_1915_ ),
    .B1(\heichips25_sap3/net76 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][1] ),
    .A2(\heichips25_sap3/net83 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][1] ));
 sg13g2_and2_1 \heichips25_sap3/_2503_  (.A(\heichips25_sap3/_1914_ ),
    .B(\heichips25_sap3/_1915_ ),
    .X(\heichips25_sap3/_1916_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_2504_  (.B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][1] ),
    .C1(\heichips25_sap3/net79 ),
    .B1(\heichips25_sap3/net78 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][1] ),
    .Y(\heichips25_sap3/_1917_ ),
    .A2(\heichips25_sap3/net218 ));
 sg13g2_a22oi_1 \heichips25_sap3/_2505_  (.Y(\heichips25_sap3/_1918_ ),
    .B1(\heichips25_sap3/net88 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][1] ),
    .A2(\heichips25_sap3/net89 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][1] ));
 sg13g2_a22oi_1 \heichips25_sap3/_2506_  (.Y(\heichips25_sap3/_1919_ ),
    .B1(\heichips25_sap3/net82 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][1] ),
    .A2(\heichips25_sap3/net86 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][1] ));
 sg13g2_and3_1 \heichips25_sap3/_2507_  (.X(\heichips25_sap3/_1920_ ),
    .A(\heichips25_sap3/_1917_ ),
    .B(\heichips25_sap3/_1918_ ),
    .C(\heichips25_sap3/_1919_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2508_  (.A1(\heichips25_sap3/_1916_ ),
    .A2(\heichips25_sap3/_1920_ ),
    .Y(\heichips25_sap3/_1921_ ),
    .B1(\heichips25_sap3/net67 ));
 sg13g2_or3_1 \heichips25_sap3/_2509_  (.A(\heichips25_sap3/_1908_ ),
    .B(\heichips25_sap3/_1913_ ),
    .C(\heichips25_sap3/_1921_ ),
    .X(\uio_out_sap3[1] ));
 sg13g2_inv_1 \heichips25_sap3/_2510_  (.Y(\heichips25_sap3/_1922_ ),
    .A(\uio_out_sap3[1] ));
 sg13g2_nor2_1 \heichips25_sap3/_2511_  (.A(\heichips25_sap3/sap_3_inst.alu_inst.carry ),
    .B(\heichips25_sap3/net215 ),
    .Y(\heichips25_sap3/_1923_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2512_  (.B1(\heichips25_sap3/_1899_ ),
    .Y(\heichips25_sap3/_1924_ ),
    .A1(\heichips25_sap3/_1802_ ),
    .A2(\uio_out_sap3[1] ));
 sg13g2_o21ai_1 \heichips25_sap3/_2513_  (.B1(\heichips25_sap3/_1900_ ),
    .Y(\heichips25_sap3/_0034_ ),
    .A1(\heichips25_sap3/_1923_ ),
    .A2(\heichips25_sap3/_1924_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2514_  (.B1(\heichips25_sap3/sap_3_inst.alu_flags[0] ),
    .Y(\heichips25_sap3/_1925_ ),
    .A1(\heichips25_sap3/_1717_ ),
    .A2(\heichips25_sap3/_1878_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2515_  (.Y(\heichips25_sap3/_1926_ ),
    .B1(\heichips25_sap3/net79 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][0] ),
    .A2(\heichips25_sap3/net86 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][0] ));
 sg13g2_a22oi_1 \heichips25_sap3/_2516_  (.Y(\heichips25_sap3/_1927_ ),
    .B1(\heichips25_sap3/net71 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][0] ),
    .A2(\heichips25_sap3/net216 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][0] ));
 sg13g2_a22oi_1 \heichips25_sap3/_2517_  (.Y(\heichips25_sap3/_1928_ ),
    .B1(\heichips25_sap3/net82 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][0] ),
    .A2(\heichips25_sap3/net88 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][0] ));
 sg13g2_a22oi_1 \heichips25_sap3/_2518_  (.Y(\heichips25_sap3/_1929_ ),
    .B1(\heichips25_sap3/net76 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][0] ),
    .A2(\heichips25_sap3/net83 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][0] ));
 sg13g2_and2_1 \heichips25_sap3/_2519_  (.A(\heichips25_sap3/_1928_ ),
    .B(\heichips25_sap3/_1929_ ),
    .X(\heichips25_sap3/_1930_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2520_  (.Y(\heichips25_sap3/_1931_ ),
    .B1(\heichips25_sap3/net74 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][0] ),
    .A2(\heichips25_sap3/net78 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][0] ));
 sg13g2_and4_1 \heichips25_sap3/_2521_  (.A(\heichips25_sap3/_1734_ ),
    .B(\heichips25_sap3/_1926_ ),
    .C(\heichips25_sap3/_1927_ ),
    .D(\heichips25_sap3/_1931_ ),
    .X(\heichips25_sap3/_0198_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_2522_  (.B2(\heichips25_sap3/_0198_ ),
    .C1(\heichips25_sap3/_1654_ ),
    .B1(\heichips25_sap3/_1930_ ),
    .A1(\heichips25_sap3/_1392_ ),
    .Y(\heichips25_sap3/_0199_ ),
    .A2(\heichips25_sap3/net89 ));
 sg13g2_and2_1 \heichips25_sap3/_2523_  (.A(net3),
    .B(\heichips25_sap3/_1770_ ),
    .X(\heichips25_sap3/_0200_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2524_  (.A(\heichips25_sap3/net289 ),
    .B(\heichips25_sap3/net156 ),
    .Y(\heichips25_sap3/_0201_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2525_  (.Y(\heichips25_sap3/_0202_ ),
    .A(\heichips25_sap3/sap_3_inst.alu_flags[0] ),
    .B(\heichips25_sap3/_1788_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2526_  (.A1(\heichips25_sap3/net156 ),
    .A2(\heichips25_sap3/_0202_ ),
    .Y(\heichips25_sap3/_0203_ ),
    .B1(\heichips25_sap3/_0201_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2527_  (.Y(\heichips25_sap3/_0204_ ),
    .B1(\heichips25_sap3/net78 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][0] ),
    .A2(\heichips25_sap3/net89 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][0] ));
 sg13g2_a22oi_1 \heichips25_sap3/_2528_  (.Y(\heichips25_sap3/_0205_ ),
    .B1(\heichips25_sap3/net74 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][0] ),
    .A2(\heichips25_sap3/net88 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][0] ));
 sg13g2_and2_1 \heichips25_sap3/_2529_  (.A(\heichips25_sap3/_0204_ ),
    .B(\heichips25_sap3/_0205_ ),
    .X(\heichips25_sap3/_0206_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2530_  (.Y(\heichips25_sap3/_0207_ ),
    .B1(\heichips25_sap3/net76 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][0] ),
    .A2(\heichips25_sap3/net83 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][0] ));
 sg13g2_a22oi_1 \heichips25_sap3/_2531_  (.Y(\heichips25_sap3/_0208_ ),
    .B1(\heichips25_sap3/net82 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][0] ),
    .A2(\heichips25_sap3/net86 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][0] ));
 sg13g2_a22oi_1 \heichips25_sap3/_2532_  (.Y(\heichips25_sap3/_0209_ ),
    .B1(\heichips25_sap3/net71 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][0] ),
    .A2(\heichips25_sap3/net216 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][0] ));
 sg13g2_and4_1 \heichips25_sap3/_2533_  (.A(\heichips25_sap3/_1742_ ),
    .B(\heichips25_sap3/_0207_ ),
    .C(\heichips25_sap3/_0208_ ),
    .D(\heichips25_sap3/_0209_ ),
    .X(\heichips25_sap3/_0210_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2534_  (.A1(\heichips25_sap3/_0206_ ),
    .A2(\heichips25_sap3/_0210_ ),
    .Y(\heichips25_sap3/_0211_ ),
    .B1(\heichips25_sap3/net67 ));
 sg13g2_or4_1 \heichips25_sap3/_2535_  (.A(\heichips25_sap3/_0199_ ),
    .B(\heichips25_sap3/_0200_ ),
    .C(\heichips25_sap3/_0203_ ),
    .D(\heichips25_sap3/_0211_ ),
    .X(\uio_out_sap3[0] ));
 sg13g2_inv_1 \heichips25_sap3/_2536_  (.Y(\heichips25_sap3/_0212_ ),
    .A(\uio_out_sap3[0] ));
 sg13g2_nor2_1 \heichips25_sap3/_2537_  (.A(\heichips25_sap3/_1883_ ),
    .B(\heichips25_sap3/_1892_ ),
    .Y(\heichips25_sap3/_0213_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2538_  (.A(\heichips25_sap3/_1886_ ),
    .B(\heichips25_sap3/_0213_ ),
    .Y(\heichips25_sap3/_0214_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2539_  (.A(\heichips25_sap3/net286 ),
    .B(\heichips25_sap3/net289 ),
    .C(\heichips25_sap3/net279 ),
    .Y(\heichips25_sap3/_0215_ ));
 sg13g2_nor4_1 \heichips25_sap3/_2540_  (.A(\heichips25_sap3/net282 ),
    .B(\heichips25_sap3/net274 ),
    .C(\heichips25_sap3/net284 ),
    .D(\heichips25_sap3/net277 ),
    .Y(\heichips25_sap3/_0216_ ));
 sg13g2_nand3_1 \heichips25_sap3/_2541_  (.B(\heichips25_sap3/_0215_ ),
    .C(\heichips25_sap3/_0216_ ),
    .A(\heichips25_sap3/_1383_ ),
    .Y(\heichips25_sap3/_0217_ ));
 sg13g2_nor4_1 \heichips25_sap3/_2542_  (.A(\heichips25_sap3/sap_3_inst.alu_inst.act[1] ),
    .B(\heichips25_sap3/sap_3_inst.alu_inst.act[0] ),
    .C(\heichips25_sap3/sap_3_inst.alu_inst.act[3] ),
    .D(\heichips25_sap3/sap_3_inst.alu_inst.act[2] ),
    .Y(\heichips25_sap3/_0218_ ));
 sg13g2_nor4_1 \heichips25_sap3/_2543_  (.A(\heichips25_sap3/sap_3_inst.alu_inst.act[5] ),
    .B(\heichips25_sap3/sap_3_inst.alu_inst.act[4] ),
    .C(\heichips25_sap3/sap_3_inst.alu_inst.act[7] ),
    .D(\heichips25_sap3/sap_3_inst.alu_inst.act[6] ),
    .Y(\heichips25_sap3/_0219_ ));
 sg13g2_nand3_1 \heichips25_sap3/_2544_  (.B(\heichips25_sap3/_0218_ ),
    .C(\heichips25_sap3/_0219_ ),
    .A(\heichips25_sap3/_0214_ ),
    .Y(\heichips25_sap3/_0220_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2545_  (.B1(\heichips25_sap3/_0220_ ),
    .Y(\heichips25_sap3/_0221_ ),
    .A1(\heichips25_sap3/_0214_ ),
    .A2(\heichips25_sap3/_0217_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2546_  (.A(\heichips25_sap3/net215 ),
    .B(\heichips25_sap3/_0221_ ),
    .Y(\heichips25_sap3/_0222_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2547_  (.A(\heichips25_sap3/_1717_ ),
    .B(\heichips25_sap3/_1878_ ),
    .C(\heichips25_sap3/_0222_ ),
    .Y(\heichips25_sap3/_0223_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2548_  (.B1(\heichips25_sap3/_0223_ ),
    .Y(\heichips25_sap3/_0224_ ),
    .A1(\heichips25_sap3/_1802_ ),
    .A2(\uio_out_sap3[0] ));
 sg13g2_nand2_1 \heichips25_sap3/_2549_  (.Y(\heichips25_sap3/_0033_ ),
    .A(\heichips25_sap3/_1925_ ),
    .B(\heichips25_sap3/_0224_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2550_  (.Y(\heichips25_sap3/_0225_ ),
    .B1(\heichips25_sap3/net73 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][3] ),
    .A2(\heichips25_sap3/net77 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][3] ));
 sg13g2_a22oi_1 \heichips25_sap3/_2551_  (.Y(\heichips25_sap3/_0226_ ),
    .B1(\heichips25_sap3/net80 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][3] ),
    .A2(\heichips25_sap3/net85 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][3] ));
 sg13g2_and2_1 \heichips25_sap3/_2552_  (.A(\heichips25_sap3/_0225_ ),
    .B(\heichips25_sap3/_0226_ ),
    .X(\heichips25_sap3/_0227_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2553_  (.Y(\heichips25_sap3/_0228_ ),
    .B1(\heichips25_sap3/net82 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][3] ),
    .A2(\heichips25_sap3/net83 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][3] ));
 sg13g2_a22oi_1 \heichips25_sap3/_2554_  (.Y(\heichips25_sap3/_0229_ ),
    .B1(\heichips25_sap3/net76 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][3] ),
    .A2(\heichips25_sap3/net216 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][3] ));
 sg13g2_a22oi_1 \heichips25_sap3/_2555_  (.Y(\heichips25_sap3/_0230_ ),
    .B1(\heichips25_sap3/net71 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][3] ),
    .A2(\heichips25_sap3/net87 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][3] ));
 sg13g2_and4_1 \heichips25_sap3/_2556_  (.A(\heichips25_sap3/_1734_ ),
    .B(\heichips25_sap3/_0228_ ),
    .C(\heichips25_sap3/_0229_ ),
    .D(\heichips25_sap3/_0230_ ),
    .X(\heichips25_sap3/_0231_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_2557_  (.B2(\heichips25_sap3/_0231_ ),
    .C1(\heichips25_sap3/_1654_ ),
    .B1(\heichips25_sap3/_0227_ ),
    .A1(\heichips25_sap3/_1368_ ),
    .Y(\heichips25_sap3/_0232_ ),
    .A2(\heichips25_sap3/net92 ));
 sg13g2_a22oi_1 \heichips25_sap3/_2558_  (.Y(\heichips25_sap3/_0233_ ),
    .B1(\heichips25_sap3/_1788_ ),
    .B2(\heichips25_sap3/sap_3_inst.alu_flags[3] ),
    .A2(\heichips25_sap3/_1770_ ),
    .A1(net6));
 sg13g2_o21ai_1 \heichips25_sap3/_2559_  (.B1(\heichips25_sap3/_0233_ ),
    .Y(\heichips25_sap3/_0234_ ),
    .A1(\heichips25_sap3/_1367_ ),
    .A2(\heichips25_sap3/net155 ));
 sg13g2_a22oi_1 \heichips25_sap3/_2560_  (.Y(\heichips25_sap3/_0235_ ),
    .B1(\heichips25_sap3/net77 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][3] ),
    .A2(\heichips25_sap3/net90 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][3] ));
 sg13g2_a22oi_1 \heichips25_sap3/_2561_  (.Y(\heichips25_sap3/_0236_ ),
    .B1(\heichips25_sap3/net75 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][3] ),
    .A2(\heichips25_sap3/net216 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][3] ));
 sg13g2_a221oi_1 \heichips25_sap3/_2562_  (.B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][3] ),
    .C1(\heichips25_sap3/net79 ),
    .B1(\heichips25_sap3/net71 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][3] ),
    .Y(\heichips25_sap3/_0237_ ),
    .A2(\heichips25_sap3/net83 ));
 sg13g2_a22oi_1 \heichips25_sap3/_2563_  (.Y(\heichips25_sap3/_0238_ ),
    .B1(\heichips25_sap3/net73 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][3] ),
    .A2(\heichips25_sap3/net81 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][3] ));
 sg13g2_a22oi_1 \heichips25_sap3/_2564_  (.Y(\heichips25_sap3/_0239_ ),
    .B1(\heichips25_sap3/net85 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][3] ),
    .A2(\heichips25_sap3/net88 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][3] ));
 sg13g2_and4_1 \heichips25_sap3/_2565_  (.A(\heichips25_sap3/_0235_ ),
    .B(\heichips25_sap3/_0236_ ),
    .C(\heichips25_sap3/_0238_ ),
    .D(\heichips25_sap3/_0239_ ),
    .X(\heichips25_sap3/_0240_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2566_  (.A1(\heichips25_sap3/_0237_ ),
    .A2(\heichips25_sap3/_0240_ ),
    .Y(\heichips25_sap3/_0241_ ),
    .B1(\heichips25_sap3/net66 ));
 sg13g2_nor3_1 \heichips25_sap3/_2567_  (.A(\heichips25_sap3/_0232_ ),
    .B(\heichips25_sap3/_0234_ ),
    .C(\heichips25_sap3/_0241_ ),
    .Y(\heichips25_sap3/_0242_ ));
 sg13g2_inv_1 \heichips25_sap3/_2568_  (.Y(\uio_out_sap3[3] ),
    .A(\heichips25_sap3/net45 ));
 sg13g2_or2_1 \heichips25_sap3/_2569_  (.X(\heichips25_sap3/_0243_ ),
    .B(\heichips25_sap3/_0214_ ),
    .A(\heichips25_sap3/_1878_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2570_  (.A1(\heichips25_sap3/net215 ),
    .A2(\heichips25_sap3/net45 ),
    .Y(\heichips25_sap3/_0244_ ),
    .B1(\heichips25_sap3/_0243_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2571_  (.B1(\heichips25_sap3/_0244_ ),
    .Y(\heichips25_sap3/_0245_ ),
    .A1(\heichips25_sap3/net275 ),
    .A2(\heichips25_sap3/_1801_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2572_  (.Y(\heichips25_sap3/_0246_ ),
    .A(\heichips25_sap3/sap_3_inst.alu_flags[3] ),
    .B(\heichips25_sap3/_0243_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2573_  (.Y(\heichips25_sap3/_0032_ ),
    .A(\heichips25_sap3/_0245_ ),
    .B(\heichips25_sap3/_0246_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2574_  (.A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[0][2] ),
    .B(\heichips25_sap3/_1734_ ),
    .Y(\heichips25_sap3/_0247_ ));
 sg13g2_nand4_1 \heichips25_sap3/_2575_  (.B(\heichips25_sap3/_1695_ ),
    .C(\heichips25_sap3/_1712_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][2] ),
    .Y(\heichips25_sap3/_0248_ ),
    .D(\heichips25_sap3/_1731_ ));
 sg13g2_nand4_1 \heichips25_sap3/_2576_  (.B(\heichips25_sap3/_1695_ ),
    .C(\heichips25_sap3/_1713_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][2] ),
    .Y(\heichips25_sap3/_0249_ ),
    .D(\heichips25_sap3/_1731_ ));
 sg13g2_nand4_1 \heichips25_sap3/_2577_  (.B(\heichips25_sap3/_1680_ ),
    .C(\heichips25_sap3/_1713_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][2] ),
    .Y(\heichips25_sap3/_0250_ ),
    .D(\heichips25_sap3/_1731_ ));
 sg13g2_nand3_1 \heichips25_sap3/_2578_  (.B(\heichips25_sap3/_1695_ ),
    .C(\heichips25_sap3/net827 ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][2] ),
    .Y(\heichips25_sap3/_0251_ ));
 sg13g2_and4_1 \heichips25_sap3/_2579_  (.A(\heichips25_sap3/_0248_ ),
    .B(\heichips25_sap3/_0249_ ),
    .C(\heichips25_sap3/_0250_ ),
    .D(\heichips25_sap3/_0251_ ),
    .X(\heichips25_sap3/_0252_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_2580_  (.B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][2] ),
    .C1(\heichips25_sap3/net89 ),
    .B1(\heichips25_sap3/net82 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][2] ),
    .Y(\heichips25_sap3/_0253_ ),
    .A2(\heichips25_sap3/net218 ));
 sg13g2_a22oi_1 \heichips25_sap3/_2581_  (.Y(\heichips25_sap3/_0254_ ),
    .B1(\heichips25_sap3/net74 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][2] ),
    .A2(\heichips25_sap3/net79 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][2] ));
 sg13g2_a22oi_1 \heichips25_sap3/_2582_  (.Y(\heichips25_sap3/_0255_ ),
    .B1(\heichips25_sap3/net76 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][2] ),
    .A2(\heichips25_sap3/net78 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][2] ));
 sg13g2_and4_1 \heichips25_sap3/_2583_  (.A(\heichips25_sap3/_0252_ ),
    .B(\heichips25_sap3/_0253_ ),
    .C(\heichips25_sap3/_0254_ ),
    .D(\heichips25_sap3/_0255_ ),
    .X(\heichips25_sap3/_0256_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2584_  (.A(\heichips25_sap3/_1654_ ),
    .B(\heichips25_sap3/_0247_ ),
    .C(\heichips25_sap3/_0256_ ),
    .Y(\heichips25_sap3/_0257_ ));
 sg13g2_and2_1 \heichips25_sap3/_2585_  (.A(net5),
    .B(\heichips25_sap3/_1770_ ),
    .X(\heichips25_sap3/_0258_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2586_  (.A(\heichips25_sap3/net284 ),
    .B(\heichips25_sap3/net156 ),
    .Y(\heichips25_sap3/_0259_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2587_  (.Y(\heichips25_sap3/_0260_ ),
    .A(\heichips25_sap3/sap_3_inst.alu_flags[2] ),
    .B(\heichips25_sap3/_1788_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2588_  (.A1(\heichips25_sap3/net156 ),
    .A2(\heichips25_sap3/_0260_ ),
    .Y(\heichips25_sap3/_0261_ ),
    .B1(\heichips25_sap3/_0259_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2589_  (.Y(\heichips25_sap3/_0262_ ),
    .B1(\heichips25_sap3/net76 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][2] ),
    .A2(\heichips25_sap3/net82 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][2] ));
 sg13g2_a22oi_1 \heichips25_sap3/_2590_  (.Y(\heichips25_sap3/_0263_ ),
    .B1(\heichips25_sap3/net78 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][2] ),
    .A2(\heichips25_sap3/net88 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][2] ));
 sg13g2_a221oi_1 \heichips25_sap3/_2591_  (.B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][2] ),
    .C1(\heichips25_sap3/net79 ),
    .B1(\heichips25_sap3/net74 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][2] ),
    .Y(\heichips25_sap3/_0264_ ),
    .A2(\heichips25_sap3/net83 ));
 sg13g2_a22oi_1 \heichips25_sap3/_2592_  (.Y(\heichips25_sap3/_0265_ ),
    .B1(\heichips25_sap3/net71 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][2] ),
    .A2(\heichips25_sap3/net218 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][2] ));
 sg13g2_a22oi_1 \heichips25_sap3/_2593_  (.Y(\heichips25_sap3/_0266_ ),
    .B1(\heichips25_sap3/net86 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][2] ),
    .A2(\heichips25_sap3/net89 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][2] ));
 sg13g2_and4_1 \heichips25_sap3/_2594_  (.A(\heichips25_sap3/_0262_ ),
    .B(\heichips25_sap3/_0263_ ),
    .C(\heichips25_sap3/_0265_ ),
    .D(\heichips25_sap3/_0266_ ),
    .X(\heichips25_sap3/_0267_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2595_  (.A1(\heichips25_sap3/_0264_ ),
    .A2(\heichips25_sap3/_0267_ ),
    .Y(\heichips25_sap3/_0268_ ),
    .B1(\heichips25_sap3/net67 ));
 sg13g2_or4_1 \heichips25_sap3/_2596_  (.A(\heichips25_sap3/_0257_ ),
    .B(\heichips25_sap3/_0258_ ),
    .C(\heichips25_sap3/_0261_ ),
    .D(\heichips25_sap3/_0268_ ),
    .X(\uio_out_sap3[2] ));
 sg13g2_nand2_1 \heichips25_sap3/_2597_  (.Y(\heichips25_sap3/_0269_ ),
    .A(\heichips25_sap3/_1801_ ),
    .B(net44));
 sg13g2_xor2_1 \heichips25_sap3/_2598_  (.B(\heichips25_sap3/net277 ),
    .A(\heichips25_sap3/net275 ),
    .X(\heichips25_sap3/_0270_ ));
 sg13g2_xor2_1 \heichips25_sap3/_2599_  (.B(\heichips25_sap3/net280 ),
    .A(\heichips25_sap3/net279 ),
    .X(\heichips25_sap3/_0271_ ));
 sg13g2_xnor2_1 \heichips25_sap3/_2600_  (.Y(\heichips25_sap3/_0272_ ),
    .A(\heichips25_sap3/_0270_ ),
    .B(\heichips25_sap3/_0271_ ));
 sg13g2_xor2_1 \heichips25_sap3/_2601_  (.B(\heichips25_sap3/net289 ),
    .A(\heichips25_sap3/net287 ),
    .X(\heichips25_sap3/_0273_ ));
 sg13g2_xor2_1 \heichips25_sap3/_2602_  (.B(\heichips25_sap3/sap_3_inst.alu_inst.acc[2] ),
    .A(\heichips25_sap3/net283 ),
    .X(\heichips25_sap3/_0274_ ));
 sg13g2_xnor2_1 \heichips25_sap3/_2603_  (.Y(\heichips25_sap3/_0275_ ),
    .A(\heichips25_sap3/_0273_ ),
    .B(\heichips25_sap3/_0274_ ));
 sg13g2_xnor2_1 \heichips25_sap3/_2604_  (.Y(\heichips25_sap3/_0276_ ),
    .A(\heichips25_sap3/_0272_ ),
    .B(\heichips25_sap3/_0275_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2605_  (.A1(\heichips25_sap3/_1802_ ),
    .A2(\heichips25_sap3/_0276_ ),
    .Y(\heichips25_sap3/_0277_ ),
    .B1(\heichips25_sap3/_0243_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2606_  (.Y(\heichips25_sap3/_0031_ ),
    .B1(\heichips25_sap3/_0269_ ),
    .B2(\heichips25_sap3/_0277_ ),
    .A2(\heichips25_sap3/_0243_ ),
    .A1(\heichips25_sap3/_1358_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_2607_  (.Y(\heichips25_sap3/_0278_ ),
    .B(\heichips25_sap3/_1636_ ),
    .A_N(\heichips25_sap3/_1553_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2608_  (.B1(\heichips25_sap3/_1635_ ),
    .Y(\heichips25_sap3/_0279_ ),
    .A1(\heichips25_sap3/_1530_ ),
    .A2(\heichips25_sap3/_1531_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2609_  (.Y(\heichips25_sap3/_0280_ ),
    .B1(\heichips25_sap3/_0279_ ),
    .B2(\heichips25_sap3/_1528_ ),
    .A2(\heichips25_sap3/_0278_ ),
    .A1(\heichips25_sap3/_1498_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_2610_  (.Y(\heichips25_sap3/_0281_ ),
    .B(\heichips25_sap3/_1514_ ),
    .A_N(\heichips25_sap3/_1561_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2611_  (.A(\heichips25_sap3/net236 ),
    .B(\heichips25_sap3/_1584_ ),
    .Y(\heichips25_sap3/_0282_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2612_  (.Y(\heichips25_sap3/_0283_ ),
    .B1(\heichips25_sap3/_0281_ ),
    .B2(\heichips25_sap3/_0282_ ),
    .A2(\heichips25_sap3/_1521_ ),
    .A1(\heichips25_sap3/_1514_ ));
 sg13g2_nand4_1 \heichips25_sap3/_2613_  (.B(\heichips25_sap3/_1484_ ),
    .C(\heichips25_sap3/_1579_ ),
    .A(\heichips25_sap3/net241 ),
    .Y(\heichips25_sap3/_0284_ ),
    .D(\heichips25_sap3/_1612_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2614_  (.A(\heichips25_sap3/_0280_ ),
    .B(\heichips25_sap3/_0283_ ),
    .C(\heichips25_sap3/_0284_ ),
    .Y(\heichips25_sap3/_0285_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2615_  (.B1(\heichips25_sap3/_1592_ ),
    .Y(\heichips25_sap3/mem_mar_we ),
    .A1(\heichips25_sap3/_1471_ ),
    .A2(\heichips25_sap3/_0285_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2616_  (.A(\heichips25_sap3/_1359_ ),
    .B(\heichips25_sap3/net1019 ),
    .Y(\heichips25_sap3/_0286_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2617_  (.Y(\heichips25_sap3/_0287_ ),
    .A(\heichips25_sap3/net1064 ),
    .B(\heichips25_sap3/_1433_ ));
 sg13g2_nor2b_1 \heichips25_sap3/_2618_  (.A(\heichips25_sap3/_0286_ ),
    .B_N(\heichips25_sap3/_0287_ ),
    .Y(\heichips25_sap3/_0288_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2619_  (.Y(\heichips25_sap3/_0001_ ),
    .A(\heichips25_sap3/_1366_ ),
    .B(\heichips25_sap3/_0288_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2620_  (.Y(\heichips25_sap3/_0289_ ),
    .A(\heichips25_sap3/net1130 ),
    .B(\heichips25_sap3/_1431_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2621_  (.A(\heichips25_sap3/_1360_ ),
    .B(\heichips25_sap3/net835 ),
    .Y(\heichips25_sap3/_0290_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2622_  (.A1(\heichips25_sap3/net1130 ),
    .A2(\heichips25_sap3/_1431_ ),
    .Y(\heichips25_sap3/_0291_ ),
    .B1(\heichips25_sap3/_0290_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_2623_  (.Y(\heichips25_sap3/_0000_ ),
    .B(\heichips25_sap3/net1131 ),
    .A_N(\heichips25_sap3/net832 ));
 sg13g2_a22oi_1 \heichips25_sap3/_2624_  (.Y(\heichips25_sap3/_0292_ ),
    .B1(\heichips25_sap3/_1682_ ),
    .B2(\heichips25_sap3/_1537_ ),
    .A2(\heichips25_sap3/_1627_ ),
    .A1(\heichips25_sap3/_1513_ ));
 sg13g2_nand4_1 \heichips25_sap3/_2625_  (.B(\heichips25_sap3/_1667_ ),
    .C(\heichips25_sap3/_1775_ ),
    .A(\heichips25_sap3/_1630_ ),
    .Y(\heichips25_sap3/_0293_ ),
    .D(\heichips25_sap3/_0292_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2626_  (.Y(\heichips25_sap3/_0294_ ),
    .B1(\heichips25_sap3/_1784_ ),
    .B2(\heichips25_sap3/_0293_ ),
    .A2(\heichips25_sap3/net228 ),
    .A1(\heichips25_sap3/net248 ));
 sg13g2_nor2_1 \heichips25_sap3/_2627_  (.A(\heichips25_sap3/_1455_ ),
    .B(\heichips25_sap3/_0294_ ),
    .Y(\heichips25_sap3/mem_ram_we ));
 sg13g2_nor4_1 \heichips25_sap3/_2628_  (.A(\heichips25_sap3/_1435_ ),
    .B(\heichips25_sap3/_1448_ ),
    .C(\heichips25_sap3/_1464_ ),
    .D(\heichips25_sap3/_1478_ ),
    .Y(\heichips25_sap3/_0295_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2629_  (.B1(\heichips25_sap3/_1559_ ),
    .Y(\heichips25_sap3/_0296_ ),
    .A1(\heichips25_sap3/_1522_ ),
    .A2(\heichips25_sap3/_1526_ ));
 sg13g2_nand4_1 \heichips25_sap3/_2630_  (.B(\heichips25_sap3/_1487_ ),
    .C(\heichips25_sap3/_1502_ ),
    .A(\heichips25_sap3/net237 ),
    .Y(\heichips25_sap3/_0297_ ),
    .D(\heichips25_sap3/_1541_ ));
 sg13g2_nand3_1 \heichips25_sap3/_2631_  (.B(\heichips25_sap3/net244 ),
    .C(\heichips25_sap3/_1551_ ),
    .A(\heichips25_sap3/_1459_ ),
    .Y(\heichips25_sap3/_0298_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2632_  (.A1(\heichips25_sap3/_1503_ ),
    .A2(\heichips25_sap3/_1568_ ),
    .Y(\heichips25_sap3/_0299_ ),
    .B1(\heichips25_sap3/_0295_ ));
 sg13g2_nand4_1 \heichips25_sap3/_2633_  (.B(\heichips25_sap3/_1718_ ),
    .C(\heichips25_sap3/_1774_ ),
    .A(\heichips25_sap3/_1573_ ),
    .Y(\heichips25_sap3/_0300_ ),
    .D(\heichips25_sap3/_0299_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2634_  (.B1(\heichips25_sap3/_1568_ ),
    .Y(\heichips25_sap3/_0301_ ),
    .A1(\heichips25_sap3/_1491_ ),
    .A2(\heichips25_sap3/_1494_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2635_  (.A1(\heichips25_sap3/_0297_ ),
    .A2(\heichips25_sap3/_0301_ ),
    .Y(\heichips25_sap3/_0302_ ),
    .B1(\heichips25_sap3/net244 ));
 sg13g2_nand4_1 \heichips25_sap3/_2636_  (.B(\heichips25_sap3/_1725_ ),
    .C(\heichips25_sap3/_0296_ ),
    .A(\heichips25_sap3/_1621_ ),
    .Y(\heichips25_sap3/_0303_ ),
    .D(\heichips25_sap3/_0298_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2637_  (.A(\heichips25_sap3/_0300_ ),
    .B(\heichips25_sap3/_0302_ ),
    .C(\heichips25_sap3/_0303_ ),
    .Y(\heichips25_sap3/_0304_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2638_  (.A1(\heichips25_sap3/net235 ),
    .A2(\heichips25_sap3/_1560_ ),
    .Y(\heichips25_sap3/_0305_ ),
    .B1(\heichips25_sap3/_1558_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2639_  (.A1(\heichips25_sap3/net235 ),
    .A2(\heichips25_sap3/_1569_ ),
    .Y(\heichips25_sap3/_0306_ ),
    .B1(\heichips25_sap3/_1565_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2640_  (.A1(\heichips25_sap3/net236 ),
    .A2(\heichips25_sap3/_1543_ ),
    .Y(\heichips25_sap3/_0307_ ),
    .B1(\heichips25_sap3/_1532_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2641_  (.B1(\heichips25_sap3/_1544_ ),
    .Y(\heichips25_sap3/_0308_ ),
    .A1(\heichips25_sap3/_0305_ ),
    .A2(\heichips25_sap3/_0306_ ));
 sg13g2_nand4_1 \heichips25_sap3/_2642_  (.B(\heichips25_sap3/_1487_ ),
    .C(\heichips25_sap3/_1502_ ),
    .A(\heichips25_sap3/net237 ),
    .Y(\heichips25_sap3/_0309_ ),
    .D(\heichips25_sap3/_1541_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2643_  (.Y(\heichips25_sap3/_0310_ ),
    .A(\heichips25_sap3/_0304_ ),
    .B(\heichips25_sap3/_0308_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2644_  (.A1(\heichips25_sap3/_1576_ ),
    .A2(\heichips25_sap3/_0307_ ),
    .Y(\heichips25_sap3/_0311_ ),
    .B1(\heichips25_sap3/_0310_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2645_  (.Y(\heichips25_sap3/_0312_ ),
    .B1(\heichips25_sap3/_1623_ ),
    .B2(\heichips25_sap3/net230 ),
    .A2(\heichips25_sap3/_1605_ ),
    .A1(\heichips25_sap3/_1476_ ));
 sg13g2_and2_1 \heichips25_sap3/_2646_  (.A(\heichips25_sap3/_1719_ ),
    .B(\heichips25_sap3/_0312_ ),
    .X(\heichips25_sap3/_0313_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2647_  (.Y(\heichips25_sap3/_0314_ ),
    .A(\heichips25_sap3/_1719_ ),
    .B(\heichips25_sap3/_0312_ ));
 sg13g2_nand3_1 \heichips25_sap3/_2648_  (.B(\heichips25_sap3/_1618_ ),
    .C(\heichips25_sap3/_1643_ ),
    .A(\heichips25_sap3/net237 ),
    .Y(\heichips25_sap3/_0315_ ));
 sg13g2_nand3_1 \heichips25_sap3/_2649_  (.B(\heichips25_sap3/net224 ),
    .C(\heichips25_sap3/_0315_ ),
    .A(\heichips25_sap3/_1480_ ),
    .Y(\heichips25_sap3/_0316_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2650_  (.B1(\heichips25_sap3/_0316_ ),
    .Y(\heichips25_sap3/_0317_ ),
    .A1(\heichips25_sap3/_1875_ ),
    .A2(\heichips25_sap3/_0314_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2651_  (.B1(\heichips25_sap3/_1641_ ),
    .Y(\heichips25_sap3/_0318_ ),
    .A1(\heichips25_sap3/_0311_ ),
    .A2(\heichips25_sap3/_0317_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2652_  (.A1(\heichips25_sap3/net238 ),
    .A2(\heichips25_sap3/_1640_ ),
    .Y(\heichips25_sap3/_0319_ ),
    .B1(\heichips25_sap3/_1784_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2653_  (.A(\heichips25_sap3/net249 ),
    .B(\heichips25_sap3/net248 ),
    .C(\heichips25_sap3/_0319_ ),
    .Y(\heichips25_sap3/_0320_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2654_  (.B1(\heichips25_sap3/net227 ),
    .Y(\heichips25_sap3/_0321_ ),
    .A1(\heichips25_sap3/net249 ),
    .A2(\heichips25_sap3/net248 ));
 sg13g2_a21oi_1 \heichips25_sap3/_2655_  (.A1(\heichips25_sap3/_0318_ ),
    .A2(\heichips25_sap3/_0320_ ),
    .Y(\heichips25_sap3/_0322_ ),
    .B1(\heichips25_sap3/_1455_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2656_  (.Y(\heichips25_sap3/_0323_ ),
    .B1(\heichips25_sap3/_0321_ ),
    .B2(\heichips25_sap3/_0322_ ),
    .A2(\heichips25_sap3/net248 ),
    .A1(\heichips25_sap3/_1447_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2657_  (.Y(\heichips25_sap3/_0324_ ),
    .A(\heichips25_sap3/_1679_ ),
    .B(\heichips25_sap3/_0323_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2658_  (.A1(\heichips25_sap3/_1679_ ),
    .A2(\heichips25_sap3/_0323_ ),
    .Y(\heichips25_sap3/_0003_ ),
    .B1(\heichips25_sap3/sap_3_inst.controller_inst.stage[0] ));
 sg13g2_and2_1 \heichips25_sap3/_2659_  (.A(\heichips25_sap3/_1468_ ),
    .B(\heichips25_sap3/_0324_ ),
    .X(\heichips25_sap3/_0004_ ));
 sg13g2_xnor2_1 \heichips25_sap3/_2660_  (.Y(\heichips25_sap3/_0325_ ),
    .A(\heichips25_sap3/sap_3_inst.controller_inst.stage[2] ),
    .B(\heichips25_sap3/_1459_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2661_  (.A(\heichips25_sap3/_0323_ ),
    .B(\heichips25_sap3/_0325_ ),
    .Y(\heichips25_sap3/_0005_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2662_  (.Y(\heichips25_sap3/_0326_ ),
    .A(\heichips25_sap3/sap_3_inst.controller_inst.stage[3] ),
    .B(\heichips25_sap3/_1554_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2663_  (.A1(\heichips25_sap3/_1606_ ),
    .A2(\heichips25_sap3/_0326_ ),
    .Y(\heichips25_sap3/_0006_ ),
    .B1(\heichips25_sap3/_0323_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_2664_  (.B2(\heichips25_sap3/_0198_ ),
    .C1(\heichips25_sap3/net67 ),
    .B1(\heichips25_sap3/_1930_ ),
    .A1(\heichips25_sap3/_1392_ ),
    .Y(\uio_oe_sap3[0] ),
    .A2(\heichips25_sap3/net92 ));
 sg13g2_a221oi_1 \heichips25_sap3/_2665_  (.B2(\heichips25_sap3/_1907_ ),
    .C1(\heichips25_sap3/net67 ),
    .B1(\heichips25_sap3/_1904_ ),
    .A1(\heichips25_sap3/_1385_ ),
    .Y(\uio_oe_sap3[1] ),
    .A2(\heichips25_sap3/net89 ));
 sg13g2_inv_1 \heichips25_sap3/_2666_  (.Y(\heichips25_sap3/_0327_ ),
    .A(\uio_oe_sap3[1] ));
 sg13g2_nor3_1 \heichips25_sap3/_2667_  (.A(\heichips25_sap3/net67 ),
    .B(\heichips25_sap3/_0247_ ),
    .C(\heichips25_sap3/_0256_ ),
    .Y(\uio_oe_sap3[2] ));
 sg13g2_a221oi_1 \heichips25_sap3/_2668_  (.B2(\heichips25_sap3/_0231_ ),
    .C1(\heichips25_sap3/net66 ),
    .B1(\heichips25_sap3/_0227_ ),
    .A1(\heichips25_sap3/_1368_ ),
    .Y(\uio_oe_sap3[3] ),
    .A2(\heichips25_sap3/net92 ));
 sg13g2_inv_1 \heichips25_sap3/_2669_  (.Y(\heichips25_sap3/_0328_ ),
    .A(\uio_oe_sap3[3] ));
 sg13g2_a221oi_1 \heichips25_sap3/_2670_  (.B2(\heichips25_sap3/_1848_ ),
    .C1(\heichips25_sap3/net66 ),
    .B1(\heichips25_sap3/_1851_ ),
    .A1(\heichips25_sap3/_1400_ ),
    .Y(\uio_oe_sap3[4] ),
    .A2(\heichips25_sap3/net90 ));
 sg13g2_a221oi_1 \heichips25_sap3/_2671_  (.B2(\heichips25_sap3/_1827_ ),
    .C1(\heichips25_sap3/net66 ),
    .B1(\heichips25_sap3/_1830_ ),
    .A1(\heichips25_sap3/_1404_ ),
    .Y(\uio_oe_sap3[5] ),
    .A2(\heichips25_sap3/net91 ));
 sg13g2_nor3_1 \heichips25_sap3/_2672_  (.A(\heichips25_sap3/_1593_ ),
    .B(\heichips25_sap3/_1803_ ),
    .C(\heichips25_sap3/_1811_ ),
    .Y(\uio_oe_sap3[6] ));
 sg13g2_a221oi_1 \heichips25_sap3/_2673_  (.B2(\heichips25_sap3/_1751_ ),
    .C1(\heichips25_sap3/_1593_ ),
    .B1(\heichips25_sap3/_1747_ ),
    .A1(\heichips25_sap3/_1420_ ),
    .Y(\uio_oe_sap3[7] ),
    .A2(\heichips25_sap3/net91 ));
 sg13g2_nand3_1 \heichips25_sap3/_2674_  (.B(\heichips25_sap3/_1451_ ),
    .C(\heichips25_sap3/net237 ),
    .A(\heichips25_sap3/_1443_ ),
    .Y(\heichips25_sap3/_0002_ ));
 sg13g2_mux2_1 \heichips25_sap3/_2675_  (.A0(\heichips25_sap3/net288 ),
    .A1(\heichips25_sap3/sap_3_inst.out[0] ),
    .S(\heichips25_sap3/_0297_ ),
    .X(\heichips25_sap3/_0023_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2676_  (.Y(\heichips25_sap3/_0329_ ),
    .A(\heichips25_sap3/sap_3_inst.out[1] ),
    .B(\heichips25_sap3/net214 ));
 sg13g2_o21ai_1 \heichips25_sap3/_2677_  (.B1(\heichips25_sap3/_0329_ ),
    .Y(\heichips25_sap3/_0024_ ),
    .A1(\heichips25_sap3/_1381_ ),
    .A2(\heichips25_sap3/net214 ));
 sg13g2_mux2_1 \heichips25_sap3/_2678_  (.A0(\heichips25_sap3/net285 ),
    .A1(\heichips25_sap3/sap_3_inst.out[2] ),
    .S(\heichips25_sap3/_0297_ ),
    .X(\heichips25_sap3/_0025_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2679_  (.Y(\heichips25_sap3/_0330_ ),
    .A(\heichips25_sap3/sap_3_inst.out[3] ),
    .B(\heichips25_sap3/net213 ));
 sg13g2_o21ai_1 \heichips25_sap3/_2680_  (.B1(\heichips25_sap3/_0330_ ),
    .Y(\heichips25_sap3/_0026_ ),
    .A1(\heichips25_sap3/_1367_ ),
    .A2(\heichips25_sap3/net213 ));
 sg13g2_nand2_1 \heichips25_sap3/_2681_  (.Y(\heichips25_sap3/_0331_ ),
    .A(\heichips25_sap3/sap_3_inst.out[4] ),
    .B(\heichips25_sap3/net213 ));
 sg13g2_o21ai_1 \heichips25_sap3/_2682_  (.B1(\heichips25_sap3/_0331_ ),
    .Y(\heichips25_sap3/_0027_ ),
    .A1(\heichips25_sap3/_1383_ ),
    .A2(\heichips25_sap3/net213 ));
 sg13g2_nand2_1 \heichips25_sap3/_2683_  (.Y(\heichips25_sap3/_0332_ ),
    .A(\heichips25_sap3/sap_3_inst.out[5] ),
    .B(\heichips25_sap3/net213 ));
 sg13g2_o21ai_1 \heichips25_sap3/_2684_  (.B1(\heichips25_sap3/_0332_ ),
    .Y(\heichips25_sap3/_0028_ ),
    .A1(\heichips25_sap3/_1382_ ),
    .A2(\heichips25_sap3/net213 ));
 sg13g2_nand2_1 \heichips25_sap3/_2685_  (.Y(\heichips25_sap3/_0333_ ),
    .A(\heichips25_sap3/sap_3_inst.out[6] ),
    .B(\heichips25_sap3/net213 ));
 sg13g2_o21ai_1 \heichips25_sap3/_2686_  (.B1(\heichips25_sap3/_0333_ ),
    .Y(\heichips25_sap3/_0029_ ),
    .A1(\heichips25_sap3/_1384_ ),
    .A2(\heichips25_sap3/net213 ));
 sg13g2_nand2_1 \heichips25_sap3/_2687_  (.Y(\heichips25_sap3/_0334_ ),
    .A(\heichips25_sap3/sap_3_inst.out[7] ),
    .B(\heichips25_sap3/net214 ));
 sg13g2_o21ai_1 \heichips25_sap3/_2688_  (.B1(\heichips25_sap3/_0334_ ),
    .Y(\heichips25_sap3/_0030_ ),
    .A1(\heichips25_sap3/_1374_ ),
    .A2(\heichips25_sap3/net214 ));
 sg13g2_nor2b_1 \heichips25_sap3/_2689_  (.A(\heichips25_sap3/_1898_ ),
    .B_N(\heichips25_sap3/_1877_ ),
    .Y(\heichips25_sap3/_0335_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_2690_  (.Y(\heichips25_sap3/_0336_ ),
    .B(\heichips25_sap3/sap_3_inst.alu_inst.carry ),
    .A_N(\heichips25_sap3/_0335_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2691_  (.Y(\heichips25_sap3/_0337_ ),
    .A(\heichips25_sap3/_1884_ ),
    .B(\heichips25_sap3/net168 ));
 sg13g2_nor2_1 \heichips25_sap3/_2692_  (.A(\heichips25_sap3/_1887_ ),
    .B(\heichips25_sap3/_0337_ ),
    .Y(\heichips25_sap3/_0338_ ));
 sg13g2_or2_1 \heichips25_sap3/_2693_  (.X(\heichips25_sap3/_0339_ ),
    .B(\heichips25_sap3/_0337_ ),
    .A(\heichips25_sap3/_1887_ ));
 sg13g2_and2_1 \heichips25_sap3/_2694_  (.A(\heichips25_sap3/_1886_ ),
    .B(\heichips25_sap3/_1892_ ),
    .X(\heichips25_sap3/_0340_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2695_  (.Y(\heichips25_sap3/_0341_ ),
    .A(\heichips25_sap3/_1886_ ),
    .B(\heichips25_sap3/_1892_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2696_  (.Y(\heichips25_sap3/_0342_ ),
    .A(\heichips25_sap3/_0339_ ),
    .B(\heichips25_sap3/_0341_ ));
 sg13g2_nor2b_1 \heichips25_sap3/_2697_  (.A(\heichips25_sap3/_1887_ ),
    .B_N(\heichips25_sap3/_1894_ ),
    .Y(\heichips25_sap3/_0343_ ));
 sg13g2_nor4_1 \heichips25_sap3/_2698_  (.A(\heichips25_sap3/_1896_ ),
    .B(\heichips25_sap3/_0213_ ),
    .C(\heichips25_sap3/_0342_ ),
    .D(\heichips25_sap3/net154 ),
    .Y(\heichips25_sap3/_0344_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2699_  (.Y(\heichips25_sap3/_0345_ ),
    .A(\heichips25_sap3/_1888_ ),
    .B(\heichips25_sap3/_0344_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2700_  (.Y(\heichips25_sap3/_0346_ ),
    .A(\heichips25_sap3/_0339_ ),
    .B(\heichips25_sap3/_0345_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2701_  (.A(\heichips25_sap3/net274 ),
    .B(\heichips25_sap3/sap_3_inst.alu_inst.tmp[7] ),
    .Y(\heichips25_sap3/_0347_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2702_  (.Y(\heichips25_sap3/_0348_ ),
    .A(\heichips25_sap3/net274 ),
    .B(\heichips25_sap3/sap_3_inst.alu_inst.tmp[7] ));
 sg13g2_nor2_1 \heichips25_sap3/_2703_  (.A(\heichips25_sap3/_1384_ ),
    .B(\heichips25_sap3/_1398_ ),
    .Y(\heichips25_sap3/_0349_ ));
 sg13g2_xor2_1 \heichips25_sap3/_2704_  (.B(\heichips25_sap3/sap_3_inst.alu_inst.tmp[6] ),
    .A(\heichips25_sap3/net276 ),
    .X(\heichips25_sap3/_0350_ ));
 sg13g2_and2_1 \heichips25_sap3/_2705_  (.A(\heichips25_sap3/net278 ),
    .B(\heichips25_sap3/sap_3_inst.alu_inst.tmp[5] ),
    .X(\heichips25_sap3/_0351_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2706_  (.Y(\heichips25_sap3/_0352_ ),
    .A(\heichips25_sap3/net278 ),
    .B(\heichips25_sap3/sap_3_inst.alu_inst.tmp[5] ));
 sg13g2_nor2_1 \heichips25_sap3/_2707_  (.A(\heichips25_sap3/net278 ),
    .B(\heichips25_sap3/sap_3_inst.alu_inst.tmp[5] ),
    .Y(\heichips25_sap3/_0353_ ));
 sg13g2_and2_1 \heichips25_sap3/_2708_  (.A(\heichips25_sap3/net280 ),
    .B(\heichips25_sap3/sap_3_inst.alu_inst.tmp[4] ),
    .X(\heichips25_sap3/_0354_ ));
 sg13g2_xnor2_1 \heichips25_sap3/_2709_  (.Y(\heichips25_sap3/_0355_ ),
    .A(\heichips25_sap3/net280 ),
    .B(\heichips25_sap3/sap_3_inst.alu_inst.tmp[4] ));
 sg13g2_inv_1 \heichips25_sap3/_2710_  (.Y(\heichips25_sap3/_0356_ ),
    .A(\heichips25_sap3/_0355_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2711_  (.Y(\heichips25_sap3/_0357_ ),
    .A(\heichips25_sap3/net282 ),
    .B(\heichips25_sap3/sap_3_inst.alu_inst.tmp[3] ));
 sg13g2_nor2_1 \heichips25_sap3/_2712_  (.A(\heichips25_sap3/net282 ),
    .B(\heichips25_sap3/sap_3_inst.alu_inst.tmp[3] ),
    .Y(\heichips25_sap3/_0358_ ));
 sg13g2_or2_1 \heichips25_sap3/_2713_  (.X(\heichips25_sap3/_0359_ ),
    .B(\heichips25_sap3/sap_3_inst.alu_inst.tmp[3] ),
    .A(\heichips25_sap3/net282 ));
 sg13g2_and2_1 \heichips25_sap3/_2714_  (.A(\heichips25_sap3/net284 ),
    .B(\heichips25_sap3/sap_3_inst.alu_inst.tmp[2] ),
    .X(\heichips25_sap3/_0360_ ));
 sg13g2_xor2_1 \heichips25_sap3/_2715_  (.B(\heichips25_sap3/sap_3_inst.alu_inst.tmp[2] ),
    .A(\heichips25_sap3/net284 ),
    .X(\heichips25_sap3/_0361_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2716_  (.A(\heichips25_sap3/_1381_ ),
    .B(\heichips25_sap3/_1396_ ),
    .Y(\heichips25_sap3/_0362_ ));
 sg13g2_xor2_1 \heichips25_sap3/_2717_  (.B(\heichips25_sap3/sap_3_inst.alu_inst.tmp[1] ),
    .A(\heichips25_sap3/net286 ),
    .X(\heichips25_sap3/_0363_ ));
 sg13g2_and2_1 \heichips25_sap3/_2718_  (.A(\heichips25_sap3/net288 ),
    .B(\heichips25_sap3/sap_3_inst.alu_inst.tmp[0] ),
    .X(\heichips25_sap3/_0364_ ));
 sg13g2_a21o_1 \heichips25_sap3/_2719_  (.A2(\heichips25_sap3/_0364_ ),
    .A1(\heichips25_sap3/_0363_ ),
    .B1(\heichips25_sap3/_0362_ ),
    .X(\heichips25_sap3/_0365_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2720_  (.A1(\heichips25_sap3/_0361_ ),
    .A2(\heichips25_sap3/_0365_ ),
    .Y(\heichips25_sap3/_0366_ ),
    .B1(\heichips25_sap3/_0360_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2721_  (.A1(\heichips25_sap3/_0357_ ),
    .A2(\heichips25_sap3/_0366_ ),
    .Y(\heichips25_sap3/_0367_ ),
    .B1(\heichips25_sap3/_0358_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2722_  (.A1(\heichips25_sap3/_0356_ ),
    .A2(\heichips25_sap3/_0367_ ),
    .Y(\heichips25_sap3/_0368_ ),
    .B1(\heichips25_sap3/_0354_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2723_  (.A1(\heichips25_sap3/_0352_ ),
    .A2(\heichips25_sap3/_0368_ ),
    .Y(\heichips25_sap3/_0369_ ),
    .B1(\heichips25_sap3/_0353_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2724_  (.A1(\heichips25_sap3/_0350_ ),
    .A2(\heichips25_sap3/_0369_ ),
    .Y(\heichips25_sap3/_0370_ ),
    .B1(\heichips25_sap3/_0349_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2725_  (.B1(\heichips25_sap3/_0348_ ),
    .Y(\heichips25_sap3/_0371_ ),
    .A1(\heichips25_sap3/_0347_ ),
    .A2(\heichips25_sap3/_0370_ ));
 sg13g2_xor2_1 \heichips25_sap3/_2726_  (.B(\heichips25_sap3/sap_3_inst.alu_inst.tmp[0] ),
    .A(\heichips25_sap3/net288 ),
    .X(\heichips25_sap3/_0372_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2727_  (.Y(\heichips25_sap3/_0373_ ),
    .A(\heichips25_sap3/net254 ),
    .B(\heichips25_sap3/_0372_ ));
 sg13g2_nand3_1 \heichips25_sap3/_2728_  (.B(\heichips25_sap3/_0363_ ),
    .C(\heichips25_sap3/_0372_ ),
    .A(\heichips25_sap3/net254 ),
    .Y(\heichips25_sap3/_0374_ ));
 sg13g2_xnor2_1 \heichips25_sap3/_2729_  (.Y(\heichips25_sap3/_0375_ ),
    .A(\heichips25_sap3/_0361_ ),
    .B(\heichips25_sap3/_0365_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2730_  (.A(\heichips25_sap3/_0374_ ),
    .B(\heichips25_sap3/_0375_ ),
    .Y(\heichips25_sap3/_0376_ ));
 sg13g2_and2_1 \heichips25_sap3/_2731_  (.A(\heichips25_sap3/_0357_ ),
    .B(\heichips25_sap3/_0359_ ),
    .X(\heichips25_sap3/_0377_ ));
 sg13g2_xor2_1 \heichips25_sap3/_2732_  (.B(\heichips25_sap3/_0377_ ),
    .A(\heichips25_sap3/_0366_ ),
    .X(\heichips25_sap3/_0378_ ));
 sg13g2_or3_1 \heichips25_sap3/_2733_  (.A(\heichips25_sap3/_0374_ ),
    .B(\heichips25_sap3/_0375_ ),
    .C(\heichips25_sap3/_0378_ ),
    .X(\heichips25_sap3/_0379_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2734_  (.A(\heichips25_sap3/_0351_ ),
    .B(\heichips25_sap3/_0353_ ),
    .Y(\heichips25_sap3/_0380_ ));
 sg13g2_nor2b_1 \heichips25_sap3/_2735_  (.A(\heichips25_sap3/_0347_ ),
    .B_N(\heichips25_sap3/_0348_ ),
    .Y(\heichips25_sap3/_0381_ ));
 sg13g2_nand3_1 \heichips25_sap3/_2736_  (.B(\heichips25_sap3/_0380_ ),
    .C(\heichips25_sap3/_0381_ ),
    .A(\heichips25_sap3/_0350_ ),
    .Y(\heichips25_sap3/_0382_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2737_  (.A(\heichips25_sap3/_0355_ ),
    .B(\heichips25_sap3/_0379_ ),
    .C(\heichips25_sap3/_0382_ ),
    .Y(\heichips25_sap3/_0383_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2738_  (.B1(\heichips25_sap3/_0346_ ),
    .Y(\heichips25_sap3/_0384_ ),
    .A1(\heichips25_sap3/_0371_ ),
    .A2(\heichips25_sap3/_0383_ ));
 sg13g2_nor2b_1 \heichips25_sap3/_2739_  (.A(\heichips25_sap3/net279 ),
    .B_N(\heichips25_sap3/sap_3_inst.alu_inst.tmp[5] ),
    .Y(\heichips25_sap3/_0385_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_2740_  (.Y(\heichips25_sap3/_0386_ ),
    .B(\heichips25_sap3/net279 ),
    .A_N(\heichips25_sap3/sap_3_inst.alu_inst.tmp[5] ));
 sg13g2_nand2b_1 \heichips25_sap3/_2741_  (.Y(\heichips25_sap3/_0387_ ),
    .B(\heichips25_sap3/net283 ),
    .A_N(\heichips25_sap3/sap_3_inst.alu_inst.tmp[3] ));
 sg13g2_nor2b_1 \heichips25_sap3/_2742_  (.A(\heichips25_sap3/net283 ),
    .B_N(\heichips25_sap3/sap_3_inst.alu_inst.tmp[3] ),
    .Y(\heichips25_sap3/_0388_ ));
 sg13g2_nor2b_1 \heichips25_sap3/_2743_  (.A(\heichips25_sap3/net288 ),
    .B_N(\heichips25_sap3/sap_3_inst.alu_inst.tmp[0] ),
    .Y(\heichips25_sap3/_0389_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2744_  (.A(\heichips25_sap3/_0363_ ),
    .B(\heichips25_sap3/_0389_ ),
    .Y(\heichips25_sap3/_0390_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2745_  (.A1(\heichips25_sap3/net286 ),
    .A2(\heichips25_sap3/_1396_ ),
    .Y(\heichips25_sap3/_0391_ ),
    .B1(\heichips25_sap3/_0390_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2746_  (.A(\heichips25_sap3/_0361_ ),
    .B(\heichips25_sap3/_0391_ ),
    .Y(\heichips25_sap3/_0392_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2747_  (.A1(\heichips25_sap3/net284 ),
    .A2(\heichips25_sap3/_1397_ ),
    .Y(\heichips25_sap3/_0393_ ),
    .B1(\heichips25_sap3/_0392_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2748_  (.A1(\heichips25_sap3/_0387_ ),
    .A2(\heichips25_sap3/_0393_ ),
    .Y(\heichips25_sap3/_0394_ ),
    .B1(\heichips25_sap3/_0388_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2749_  (.A(\heichips25_sap3/_1383_ ),
    .B(\heichips25_sap3/sap_3_inst.alu_inst.tmp[4] ),
    .Y(\heichips25_sap3/_0395_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2750_  (.A1(\heichips25_sap3/_0355_ ),
    .A2(\heichips25_sap3/_0394_ ),
    .Y(\heichips25_sap3/_0396_ ),
    .B1(\heichips25_sap3/_0395_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2751_  (.B1(\heichips25_sap3/_0386_ ),
    .Y(\heichips25_sap3/_0397_ ),
    .A1(\heichips25_sap3/_0385_ ),
    .A2(\heichips25_sap3/_0396_ ));
 sg13g2_nor2b_1 \heichips25_sap3/_2752_  (.A(\heichips25_sap3/_0350_ ),
    .B_N(\heichips25_sap3/_0397_ ),
    .Y(\heichips25_sap3/_0398_ ));
 sg13g2_xnor2_1 \heichips25_sap3/_2753_  (.Y(\heichips25_sap3/_0399_ ),
    .A(\heichips25_sap3/_0350_ ),
    .B(\heichips25_sap3/_0397_ ));
 sg13g2_xor2_1 \heichips25_sap3/_2754_  (.B(\heichips25_sap3/_0389_ ),
    .A(\heichips25_sap3/_0363_ ),
    .X(\heichips25_sap3/_0400_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_2755_  (.Y(\heichips25_sap3/_0401_ ),
    .B(\heichips25_sap3/sap_3_inst.alu_flags[1] ),
    .A_N(\heichips25_sap3/_0372_ ));
 sg13g2_or2_1 \heichips25_sap3/_2756_  (.X(\heichips25_sap3/_0402_ ),
    .B(\heichips25_sap3/_0401_ ),
    .A(\heichips25_sap3/_0400_ ));
 sg13g2_xor2_1 \heichips25_sap3/_2757_  (.B(\heichips25_sap3/_0391_ ),
    .A(\heichips25_sap3/_0361_ ),
    .X(\heichips25_sap3/_0403_ ));
 sg13g2_xor2_1 \heichips25_sap3/_2758_  (.B(\heichips25_sap3/_0393_ ),
    .A(\heichips25_sap3/_0377_ ),
    .X(\heichips25_sap3/_0404_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2759_  (.A(\heichips25_sap3/_0361_ ),
    .B(\heichips25_sap3/_0377_ ),
    .C(\heichips25_sap3/_0402_ ),
    .Y(\heichips25_sap3/_0405_ ));
 sg13g2_xnor2_1 \heichips25_sap3/_2760_  (.Y(\heichips25_sap3/_0406_ ),
    .A(\heichips25_sap3/_0356_ ),
    .B(\heichips25_sap3/_0394_ ));
 sg13g2_nor2b_1 \heichips25_sap3/_2761_  (.A(\heichips25_sap3/_0406_ ),
    .B_N(\heichips25_sap3/_0405_ ),
    .Y(\heichips25_sap3/_0407_ ));
 sg13g2_xnor2_1 \heichips25_sap3/_2762_  (.Y(\heichips25_sap3/_0408_ ),
    .A(\heichips25_sap3/_0380_ ),
    .B(\heichips25_sap3/_0396_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2763_  (.Y(\heichips25_sap3/_0409_ ),
    .A(\heichips25_sap3/_0407_ ),
    .B(\heichips25_sap3/_0408_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2764_  (.A(\heichips25_sap3/_0399_ ),
    .B(\heichips25_sap3/_0409_ ),
    .Y(\heichips25_sap3/_0410_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2765_  (.A1(\heichips25_sap3/net276 ),
    .A2(\heichips25_sap3/_1398_ ),
    .Y(\heichips25_sap3/_0411_ ),
    .B1(\heichips25_sap3/_0398_ ));
 sg13g2_xor2_1 \heichips25_sap3/_2766_  (.B(\heichips25_sap3/_0411_ ),
    .A(\heichips25_sap3/_0381_ ),
    .X(\heichips25_sap3/_0412_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2767_  (.A(\heichips25_sap3/_0399_ ),
    .B(\heichips25_sap3/_0409_ ),
    .C(\heichips25_sap3/_0412_ ),
    .Y(\heichips25_sap3/_0413_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2768_  (.A1(\heichips25_sap3/_1374_ ),
    .A2(\heichips25_sap3/sap_3_inst.alu_inst.tmp[7] ),
    .Y(\heichips25_sap3/_0414_ ),
    .B1(\heichips25_sap3/_0411_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2769_  (.A1(\heichips25_sap3/net274 ),
    .A2(\heichips25_sap3/_1399_ ),
    .Y(\heichips25_sap3/_0415_ ),
    .B1(\heichips25_sap3/_0414_ ));
 sg13g2_and2_1 \heichips25_sap3/_2770_  (.A(\heichips25_sap3/net169 ),
    .B(\heichips25_sap3/_1896_ ),
    .X(\heichips25_sap3/_0416_ ));
 sg13g2_nor2b_1 \heichips25_sap3/_2771_  (.A(\heichips25_sap3/net169 ),
    .B_N(\heichips25_sap3/_1896_ ),
    .Y(\heichips25_sap3/_0417_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2772_  (.B1(\heichips25_sap3/_0340_ ),
    .Y(\heichips25_sap3/_0418_ ),
    .A1(\heichips25_sap3/_0413_ ),
    .A2(\heichips25_sap3/_0415_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2773_  (.Y(\heichips25_sap3/_0419_ ),
    .A(\heichips25_sap3/net154 ),
    .B(\heichips25_sap3/_0415_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2774_  (.A1(\heichips25_sap3/net254 ),
    .A2(\heichips25_sap3/net168 ),
    .Y(\heichips25_sap3/_0420_ ),
    .B1(\heichips25_sap3/_1888_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2775_  (.Y(\heichips25_sap3/_0421_ ),
    .B1(\heichips25_sap3/_0417_ ),
    .B2(\heichips25_sap3/net274 ),
    .A2(\heichips25_sap3/_0416_ ),
    .A1(\heichips25_sap3/net288 ));
 sg13g2_nand4_1 \heichips25_sap3/_2776_  (.B(\heichips25_sap3/_0418_ ),
    .C(\heichips25_sap3/_0419_ ),
    .A(\heichips25_sap3/_0384_ ),
    .Y(\heichips25_sap3/_0422_ ),
    .D(\heichips25_sap3/_0421_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2777_  (.A1(\heichips25_sap3/_1880_ ),
    .A2(\heichips25_sap3/_0420_ ),
    .Y(\heichips25_sap3/_0423_ ),
    .B1(\heichips25_sap3/_0422_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2778_  (.B1(\heichips25_sap3/_0335_ ),
    .Y(\heichips25_sap3/_0424_ ),
    .A1(\heichips25_sap3/_0345_ ),
    .A2(\heichips25_sap3/_0371_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2779_  (.B1(\heichips25_sap3/_0336_ ),
    .Y(\heichips25_sap3/_0039_ ),
    .A1(\heichips25_sap3/_0423_ ),
    .A2(\heichips25_sap3/_0424_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2780_  (.B1(\heichips25_sap3/_1518_ ),
    .Y(\heichips25_sap3/_0425_ ),
    .A1(\heichips25_sap3/_1442_ ),
    .A2(\heichips25_sap3/_1495_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2781_  (.A(\heichips25_sap3/net223 ),
    .B(\heichips25_sap3/_1727_ ),
    .Y(\heichips25_sap3/_0426_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2782_  (.Y(\heichips25_sap3/_0427_ ),
    .B1(\heichips25_sap3/_0425_ ),
    .B2(\heichips25_sap3/_1605_ ),
    .A2(\heichips25_sap3/_1762_ ),
    .A1(\heichips25_sap3/_1643_ ));
 sg13g2_nand4_1 \heichips25_sap3/_2783_  (.B(\heichips25_sap3/_1761_ ),
    .C(\heichips25_sap3/_0426_ ),
    .A(\heichips25_sap3/_1755_ ),
    .Y(\heichips25_sap3/_0428_ ),
    .D(\heichips25_sap3/_0427_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2784_  (.A1(\heichips25_sap3/_1646_ ),
    .A2(\heichips25_sap3/_0428_ ),
    .Y(\heichips25_sap3/_0429_ ),
    .B1(\heichips25_sap3/net221 ));
 sg13g2_nand3_1 \heichips25_sap3/_2785_  (.B(\heichips25_sap3/net238 ),
    .C(\heichips25_sap3/_1643_ ),
    .A(\heichips25_sap3/_1449_ ),
    .Y(\heichips25_sap3/_0430_ ));
 sg13g2_nand3_1 \heichips25_sap3/_2786_  (.B(\heichips25_sap3/_1767_ ),
    .C(\heichips25_sap3/_0430_ ),
    .A(\heichips25_sap3/net221 ),
    .Y(\heichips25_sap3/_0431_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2787_  (.Y(\heichips25_sap3/_0432_ ),
    .A(\heichips25_sap3/_1452_ ),
    .B(\heichips25_sap3/_0431_ ));
 sg13g2_nand3_1 \heichips25_sap3/_2788_  (.B(\heichips25_sap3/net228 ),
    .C(\heichips25_sap3/_1643_ ),
    .A(\heichips25_sap3/_1451_ ),
    .Y(\heichips25_sap3/_0433_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2789_  (.B1(\heichips25_sap3/_0433_ ),
    .Y(\heichips25_sap3/_0434_ ),
    .A1(\heichips25_sap3/_0429_ ),
    .A2(\heichips25_sap3/_0432_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2790_  (.B1(\heichips25_sap3/_1641_ ),
    .Y(\heichips25_sap3/_0435_ ),
    .A1(\heichips25_sap3/_1621_ ),
    .A2(\heichips25_sap3/_1773_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2791_  (.B1(\heichips25_sap3/_1783_ ),
    .Y(\heichips25_sap3/_0436_ ),
    .A1(\heichips25_sap3/_1776_ ),
    .A2(\heichips25_sap3/_0435_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2792_  (.A(\heichips25_sap3/_1877_ ),
    .B(\heichips25_sap3/net158 ),
    .C(\heichips25_sap3/net204 ),
    .Y(\heichips25_sap3/_0437_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2793_  (.A(\heichips25_sap3/_1721_ ),
    .B(\heichips25_sap3/_1886_ ),
    .Y(\heichips25_sap3/_0438_ ));
 sg13g2_nand3_1 \heichips25_sap3/_2794_  (.B(\heichips25_sap3/_1897_ ),
    .C(\heichips25_sap3/_0438_ ),
    .A(\heichips25_sap3/_1885_ ),
    .Y(\heichips25_sap3/_0439_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_2795_  (.Y(\heichips25_sap3/_0440_ ),
    .B(\heichips25_sap3/_0439_ ),
    .A_N(\heichips25_sap3/_0437_ ));
 sg13g2_nand4_1 \heichips25_sap3/_2796_  (.B(\heichips25_sap3/_1881_ ),
    .C(\heichips25_sap3/_1884_ ),
    .A(\heichips25_sap3/_1880_ ),
    .Y(\heichips25_sap3/_0441_ ),
    .D(\heichips25_sap3/net168 ));
 sg13g2_and4_1 \heichips25_sap3/_2797_  (.A(\heichips25_sap3/_1880_ ),
    .B(\heichips25_sap3/_1881_ ),
    .C(\heichips25_sap3/_1884_ ),
    .D(\heichips25_sap3/net168 ),
    .X(\heichips25_sap3/_0442_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2798_  (.A(\heichips25_sap3/_1870_ ),
    .B(\heichips25_sap3/_0442_ ),
    .Y(\heichips25_sap3/_0443_ ));
 sg13g2_and2_1 \heichips25_sap3/_2799_  (.A(\heichips25_sap3/_0344_ ),
    .B(\heichips25_sap3/_0443_ ),
    .X(\heichips25_sap3/_0444_ ));
 sg13g2_nor2b_1 \heichips25_sap3/_2800_  (.A(\heichips25_sap3/_1885_ ),
    .B_N(\heichips25_sap3/net169 ),
    .Y(\heichips25_sap3/_0445_ ));
 sg13g2_or3_1 \heichips25_sap3/_2801_  (.A(\heichips25_sap3/net154 ),
    .B(\heichips25_sap3/net64 ),
    .C(\heichips25_sap3/_0445_ ),
    .X(\heichips25_sap3/_0446_ ));
 sg13g2_or2_1 \heichips25_sap3/_2802_  (.X(\heichips25_sap3/_0447_ ),
    .B(\heichips25_sap3/_0443_ ),
    .A(\heichips25_sap3/net288 ));
 sg13g2_xor2_1 \heichips25_sap3/_2803_  (.B(\heichips25_sap3/_0372_ ),
    .A(\heichips25_sap3/net254 ),
    .X(\heichips25_sap3/_0448_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2804_  (.A(\heichips25_sap3/_1885_ ),
    .B(\heichips25_sap3/net169 ),
    .Y(\heichips25_sap3/_0449_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2805_  (.B1(\heichips25_sap3/net159 ),
    .Y(\heichips25_sap3/_0450_ ),
    .A1(\heichips25_sap3/net288 ),
    .A2(\heichips25_sap3/sap_3_inst.alu_inst.tmp[0] ));
 sg13g2_nand3_1 \heichips25_sap3/_2806_  (.B(\heichips25_sap3/_1894_ ),
    .C(\heichips25_sap3/_1896_ ),
    .A(\heichips25_sap3/net254 ),
    .Y(\heichips25_sap3/_0451_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2807_  (.Y(\heichips25_sap3/_0452_ ),
    .B1(\heichips25_sap3/_0449_ ),
    .B2(\heichips25_sap3/_0364_ ),
    .A2(\heichips25_sap3/_0416_ ),
    .A1(\heichips25_sap3/net287 ));
 sg13g2_nand4_1 \heichips25_sap3/_2808_  (.B(\heichips25_sap3/_0450_ ),
    .C(\heichips25_sap3/_0451_ ),
    .A(\heichips25_sap3/_0447_ ),
    .Y(\heichips25_sap3/_0453_ ),
    .D(\heichips25_sap3/_0452_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_2809_  (.B2(\heichips25_sap3/_0342_ ),
    .C1(\heichips25_sap3/_0453_ ),
    .B1(\heichips25_sap3/_0448_ ),
    .A1(\heichips25_sap3/_0372_ ),
    .Y(\heichips25_sap3/_0454_ ),
    .A2(\heichips25_sap3/_0446_ ));
 sg13g2_or2_1 \heichips25_sap3/_2810_  (.X(\heichips25_sap3/_0455_ ),
    .B(\heichips25_sap3/_0454_ ),
    .A(\heichips25_sap3/net204 ));
 sg13g2_a21oi_1 \heichips25_sap3/_2811_  (.A1(\heichips25_sap3/sap_3_inst.alu_inst.act[0] ),
    .A2(\heichips25_sap3/net204 ),
    .Y(\heichips25_sap3/_0456_ ),
    .B1(\heichips25_sap3/net158 ));
 sg13g2_a221oi_1 \heichips25_sap3/_2812_  (.B2(\heichips25_sap3/_0456_ ),
    .C1(\heichips25_sap3/net70 ),
    .B1(\heichips25_sap3/_0455_ ),
    .A1(\heichips25_sap3/_0212_ ),
    .Y(\heichips25_sap3/_0457_ ),
    .A2(\heichips25_sap3/net158 ));
 sg13g2_a21o_1 \heichips25_sap3/_2813_  (.A2(\heichips25_sap3/net70 ),
    .A1(\heichips25_sap3/net289 ),
    .B1(\heichips25_sap3/_0457_ ),
    .X(\heichips25_sap3/_0040_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2814_  (.B1(\heichips25_sap3/net159 ),
    .Y(\heichips25_sap3/_0458_ ),
    .A1(\heichips25_sap3/net286 ),
    .A2(\heichips25_sap3/sap_3_inst.alu_inst.tmp[1] ));
 sg13g2_o21ai_1 \heichips25_sap3/_2815_  (.B1(\heichips25_sap3/_0458_ ),
    .Y(\heichips25_sap3/_0459_ ),
    .A1(\heichips25_sap3/net286 ),
    .A2(\heichips25_sap3/_0441_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2816_  (.A1(\heichips25_sap3/net154 ),
    .A2(\heichips25_sap3/_0400_ ),
    .Y(\heichips25_sap3/_0460_ ),
    .B1(\heichips25_sap3/_0459_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2817_  (.A(\heichips25_sap3/_1381_ ),
    .B(\heichips25_sap3/_1619_ ),
    .C(\heichips25_sap3/_1714_ ),
    .Y(\heichips25_sap3/_0461_ ));
 sg13g2_xnor2_1 \heichips25_sap3/_2818_  (.Y(\heichips25_sap3/_0462_ ),
    .A(\heichips25_sap3/_1381_ ),
    .B(\heichips25_sap3/net212 ));
 sg13g2_o21ai_1 \heichips25_sap3/_2819_  (.B1(\heichips25_sap3/_1870_ ),
    .Y(\heichips25_sap3/_0463_ ),
    .A1(\heichips25_sap3/net288 ),
    .A2(\heichips25_sap3/_0462_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2820_  (.A1(\heichips25_sap3/net289 ),
    .A2(\heichips25_sap3/_0462_ ),
    .Y(\heichips25_sap3/_0464_ ),
    .B1(\heichips25_sap3/_0463_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_2821_  (.B2(\heichips25_sap3/net289 ),
    .C1(\heichips25_sap3/_0464_ ),
    .B1(\heichips25_sap3/_0417_ ),
    .A1(\heichips25_sap3/net285 ),
    .Y(\heichips25_sap3/_0465_ ),
    .A2(\heichips25_sap3/_0416_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2822_  (.Y(\heichips25_sap3/_0466_ ),
    .B1(\heichips25_sap3/_0449_ ),
    .B2(\heichips25_sap3/_0362_ ),
    .A2(\heichips25_sap3/_0445_ ),
    .A1(\heichips25_sap3/_0363_ ));
 sg13g2_xnor2_1 \heichips25_sap3/_2823_  (.Y(\heichips25_sap3/_0467_ ),
    .A(\heichips25_sap3/_0400_ ),
    .B(\heichips25_sap3/_0401_ ));
 sg13g2_xnor2_1 \heichips25_sap3/_2824_  (.Y(\heichips25_sap3/_0468_ ),
    .A(\heichips25_sap3/_0363_ ),
    .B(\heichips25_sap3/_0364_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2825_  (.A1(\heichips25_sap3/_0373_ ),
    .A2(\heichips25_sap3/_0468_ ),
    .Y(\heichips25_sap3/_0469_ ),
    .B1(\heichips25_sap3/_0339_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2826_  (.Y(\heichips25_sap3/_0470_ ),
    .B1(\heichips25_sap3/_0469_ ),
    .B2(\heichips25_sap3/_0374_ ),
    .A2(\heichips25_sap3/_0467_ ),
    .A1(\heichips25_sap3/_0340_ ));
 sg13g2_nand4_1 \heichips25_sap3/_2827_  (.B(\heichips25_sap3/_0465_ ),
    .C(\heichips25_sap3/_0466_ ),
    .A(\heichips25_sap3/_0460_ ),
    .Y(\heichips25_sap3/_0471_ ),
    .D(\heichips25_sap3/_0470_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2828_  (.A1(\heichips25_sap3/net64 ),
    .A2(\heichips25_sap3/_0468_ ),
    .Y(\heichips25_sap3/_0472_ ),
    .B1(\heichips25_sap3/net204 ));
 sg13g2_o21ai_1 \heichips25_sap3/_2829_  (.B1(\heichips25_sap3/_0472_ ),
    .Y(\heichips25_sap3/_0473_ ),
    .A1(\heichips25_sap3/net64 ),
    .A2(\heichips25_sap3/_0471_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2830_  (.A1(\heichips25_sap3/sap_3_inst.alu_inst.act[1] ),
    .A2(\heichips25_sap3/net204 ),
    .Y(\heichips25_sap3/_0474_ ),
    .B1(\heichips25_sap3/net158 ));
 sg13g2_a221oi_1 \heichips25_sap3/_2831_  (.B2(\heichips25_sap3/_0474_ ),
    .C1(\heichips25_sap3/net70 ),
    .B1(\heichips25_sap3/_0473_ ),
    .A1(\heichips25_sap3/_1922_ ),
    .Y(\heichips25_sap3/_0475_ ),
    .A2(\heichips25_sap3/net158 ));
 sg13g2_a21o_1 \heichips25_sap3/_2832_  (.A2(\heichips25_sap3/net70 ),
    .A1(\heichips25_sap3/net287 ),
    .B1(\heichips25_sap3/_0475_ ),
    .X(\heichips25_sap3/_0041_ ));
 sg13g2_nor2b_1 \heichips25_sap3/_2833_  (.A(net44),
    .B_N(\heichips25_sap3/net158 ),
    .Y(\heichips25_sap3/_0476_ ));
 sg13g2_and2_1 \heichips25_sap3/_2834_  (.A(\heichips25_sap3/_0360_ ),
    .B(\heichips25_sap3/_0449_ ),
    .X(\heichips25_sap3/_0477_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2835_  (.B1(\heichips25_sap3/net159 ),
    .Y(\heichips25_sap3/_0478_ ),
    .A1(\heichips25_sap3/net284 ),
    .A2(\heichips25_sap3/sap_3_inst.alu_inst.tmp[2] ));
 sg13g2_o21ai_1 \heichips25_sap3/_2836_  (.B1(\heichips25_sap3/_0478_ ),
    .Y(\heichips25_sap3/_0479_ ),
    .A1(\heichips25_sap3/net284 ),
    .A2(\heichips25_sap3/_0441_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2837_  (.Y(\heichips25_sap3/_0480_ ),
    .A(\heichips25_sap3/_0361_ ),
    .B(\heichips25_sap3/_0445_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2838_  (.Y(\heichips25_sap3/_0481_ ),
    .B1(\heichips25_sap3/_0417_ ),
    .B2(\heichips25_sap3/net287 ),
    .A2(\heichips25_sap3/_0416_ ),
    .A1(\heichips25_sap3/net282 ));
 sg13g2_nand2_1 \heichips25_sap3/_2839_  (.Y(\heichips25_sap3/_0482_ ),
    .A(\heichips25_sap3/net285 ),
    .B(\heichips25_sap3/net212 ));
 sg13g2_xnor2_1 \heichips25_sap3/_2840_  (.Y(\heichips25_sap3/_0483_ ),
    .A(\heichips25_sap3/net285 ),
    .B(\heichips25_sap3/net212 ));
 sg13g2_a21oi_1 \heichips25_sap3/_2841_  (.A1(\heichips25_sap3/net289 ),
    .A2(\heichips25_sap3/_0462_ ),
    .Y(\heichips25_sap3/_0484_ ),
    .B1(\heichips25_sap3/_0461_ ));
 sg13g2_and2_1 \heichips25_sap3/_2842_  (.A(\heichips25_sap3/_0483_ ),
    .B(\heichips25_sap3/_0484_ ),
    .X(\heichips25_sap3/_0485_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2843_  (.A(\heichips25_sap3/_0483_ ),
    .B(\heichips25_sap3/_0484_ ),
    .Y(\heichips25_sap3/_0486_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2844_  (.A(\heichips25_sap3/_1869_ ),
    .B(\heichips25_sap3/_0485_ ),
    .C(\heichips25_sap3/_0486_ ),
    .Y(\heichips25_sap3/_0487_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2845_  (.A1(\heichips25_sap3/net154 ),
    .A2(\heichips25_sap3/_0403_ ),
    .Y(\heichips25_sap3/_0488_ ),
    .B1(\heichips25_sap3/_0487_ ));
 sg13g2_xor2_1 \heichips25_sap3/_2846_  (.B(\heichips25_sap3/_0375_ ),
    .A(\heichips25_sap3/_0374_ ),
    .X(\heichips25_sap3/_0489_ ));
 sg13g2_xnor2_1 \heichips25_sap3/_2847_  (.Y(\heichips25_sap3/_0490_ ),
    .A(\heichips25_sap3/_0402_ ),
    .B(\heichips25_sap3/_0403_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2848_  (.Y(\heichips25_sap3/_0491_ ),
    .B1(\heichips25_sap3/_0490_ ),
    .B2(\heichips25_sap3/_0340_ ),
    .A2(\heichips25_sap3/_0489_ ),
    .A1(\heichips25_sap3/_0338_ ));
 sg13g2_nand4_1 \heichips25_sap3/_2849_  (.B(\heichips25_sap3/_0481_ ),
    .C(\heichips25_sap3/_0488_ ),
    .A(\heichips25_sap3/_0480_ ),
    .Y(\heichips25_sap3/_0492_ ),
    .D(\heichips25_sap3/_0491_ ));
 sg13g2_or4_1 \heichips25_sap3/_2850_  (.A(\heichips25_sap3/net64 ),
    .B(\heichips25_sap3/_0477_ ),
    .C(\heichips25_sap3/_0479_ ),
    .D(\heichips25_sap3/_0492_ ),
    .X(\heichips25_sap3/_0493_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2851_  (.A1(\heichips25_sap3/_0375_ ),
    .A2(\heichips25_sap3/net64 ),
    .Y(\heichips25_sap3/_0494_ ),
    .B1(\heichips25_sap3/net204 ));
 sg13g2_a221oi_1 \heichips25_sap3/_2852_  (.B2(\heichips25_sap3/_0494_ ),
    .C1(\heichips25_sap3/net158 ),
    .B1(\heichips25_sap3/_0493_ ),
    .A1(\heichips25_sap3/sap_3_inst.alu_inst.act[2] ),
    .Y(\heichips25_sap3/_0495_ ),
    .A2(\heichips25_sap3/net204 ));
 sg13g2_nor3_1 \heichips25_sap3/_2853_  (.A(\heichips25_sap3/net70 ),
    .B(\heichips25_sap3/_0476_ ),
    .C(\heichips25_sap3/_0495_ ),
    .Y(\heichips25_sap3/_0496_ ));
 sg13g2_a21o_1 \heichips25_sap3/_2854_  (.A2(\heichips25_sap3/net70 ),
    .A1(\heichips25_sap3/net285 ),
    .B1(\heichips25_sap3/_0496_ ),
    .X(\heichips25_sap3/_0042_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2855_  (.B1(\heichips25_sap3/_0404_ ),
    .Y(\heichips25_sap3/_0497_ ),
    .A1(\heichips25_sap3/_0402_ ),
    .A2(\heichips25_sap3/_0403_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_2856_  (.Y(\heichips25_sap3/_0498_ ),
    .B(\heichips25_sap3/_0497_ ),
    .A_N(\heichips25_sap3/_0405_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_2857_  (.Y(\heichips25_sap3/_0499_ ),
    .B(\heichips25_sap3/_0449_ ),
    .A_N(\heichips25_sap3/_0357_ ));
 sg13g2_xnor2_1 \heichips25_sap3/_2858_  (.Y(\heichips25_sap3/_0500_ ),
    .A(\heichips25_sap3/_0376_ ),
    .B(\heichips25_sap3/_0378_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2859_  (.A(\heichips25_sap3/_1367_ ),
    .B(\heichips25_sap3/_1619_ ),
    .C(\heichips25_sap3/_1714_ ),
    .Y(\heichips25_sap3/_0501_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2860_  (.A1(\heichips25_sap3/net285 ),
    .A2(\heichips25_sap3/net211 ),
    .Y(\heichips25_sap3/_0502_ ),
    .B1(\heichips25_sap3/_0486_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2861_  (.B1(\heichips25_sap3/_0482_ ),
    .Y(\heichips25_sap3/_0503_ ),
    .A1(\heichips25_sap3/_0483_ ),
    .A2(\heichips25_sap3/_0484_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2862_  (.B1(\heichips25_sap3/_1367_ ),
    .Y(\heichips25_sap3/_0504_ ),
    .A1(\heichips25_sap3/_1619_ ),
    .A2(\heichips25_sap3/_1714_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_2863_  (.Y(\heichips25_sap3/_0505_ ),
    .B(\heichips25_sap3/_0504_ ),
    .A_N(\heichips25_sap3/_0501_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2864_  (.A1(\heichips25_sap3/_0502_ ),
    .A2(\heichips25_sap3/_0505_ ),
    .Y(\heichips25_sap3/_0506_ ),
    .B1(\heichips25_sap3/_1869_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2865_  (.B1(\heichips25_sap3/_0506_ ),
    .Y(\heichips25_sap3/_0507_ ),
    .A1(\heichips25_sap3/_0502_ ),
    .A2(\heichips25_sap3/_0505_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2866_  (.Y(\heichips25_sap3/_0508_ ),
    .B1(\heichips25_sap3/_0500_ ),
    .B2(\heichips25_sap3/_0338_ ),
    .A2(\heichips25_sap3/_0498_ ),
    .A1(\heichips25_sap3/_0340_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2867_  (.Y(\heichips25_sap3/_0509_ ),
    .B1(\heichips25_sap3/_0445_ ),
    .B2(\heichips25_sap3/_0377_ ),
    .A2(\heichips25_sap3/_0404_ ),
    .A1(\heichips25_sap3/net154 ));
 sg13g2_a22oi_1 \heichips25_sap3/_2868_  (.Y(\heichips25_sap3/_0510_ ),
    .B1(\heichips25_sap3/_0417_ ),
    .B2(\heichips25_sap3/net285 ),
    .A2(\heichips25_sap3/_0359_ ),
    .A1(\heichips25_sap3/net159 ));
 sg13g2_and4_1 \heichips25_sap3/_2869_  (.A(\heichips25_sap3/_0499_ ),
    .B(\heichips25_sap3/_0508_ ),
    .C(\heichips25_sap3/_0509_ ),
    .D(\heichips25_sap3/_0510_ ),
    .X(\heichips25_sap3/_0511_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2870_  (.Y(\heichips25_sap3/_0512_ ),
    .B1(\heichips25_sap3/_0442_ ),
    .B2(\heichips25_sap3/_1367_ ),
    .A2(\heichips25_sap3/_0416_ ),
    .A1(\heichips25_sap3/net280 ));
 sg13g2_nand3_1 \heichips25_sap3/_2871_  (.B(\heichips25_sap3/_0511_ ),
    .C(\heichips25_sap3/_0512_ ),
    .A(\heichips25_sap3/_0507_ ),
    .Y(\heichips25_sap3/_0513_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2872_  (.A1(\heichips25_sap3/_0378_ ),
    .A2(\heichips25_sap3/net64 ),
    .Y(\heichips25_sap3/_0514_ ),
    .B1(\heichips25_sap3/net203 ));
 sg13g2_o21ai_1 \heichips25_sap3/_2873_  (.B1(\heichips25_sap3/_0514_ ),
    .Y(\heichips25_sap3/_0515_ ),
    .A1(\heichips25_sap3/net64 ),
    .A2(\heichips25_sap3/_0513_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2874_  (.A1(\heichips25_sap3/sap_3_inst.alu_inst.act[3] ),
    .A2(\heichips25_sap3/net203 ),
    .Y(\heichips25_sap3/_0516_ ),
    .B1(\heichips25_sap3/net157 ));
 sg13g2_a221oi_1 \heichips25_sap3/_2875_  (.B2(\heichips25_sap3/_0516_ ),
    .C1(\heichips25_sap3/net69 ),
    .B1(\heichips25_sap3/_0515_ ),
    .A1(\heichips25_sap3/net45 ),
    .Y(\heichips25_sap3/_0517_ ),
    .A2(\heichips25_sap3/net157 ));
 sg13g2_a21o_1 \heichips25_sap3/_2876_  (.A2(\heichips25_sap3/net69 ),
    .A1(\heichips25_sap3/net283 ),
    .B1(\heichips25_sap3/_0517_ ),
    .X(\heichips25_sap3/_0043_ ));
 sg13g2_nor2b_1 \heichips25_sap3/_2877_  (.A(net46),
    .B_N(\heichips25_sap3/net157 ),
    .Y(\heichips25_sap3/_0518_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2878_  (.Y(\heichips25_sap3/_0519_ ),
    .A(\heichips25_sap3/_0354_ ),
    .B(\heichips25_sap3/_0449_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2879_  (.B1(\heichips25_sap3/net159 ),
    .Y(\heichips25_sap3/_0520_ ),
    .A1(\heichips25_sap3/net281 ),
    .A2(\heichips25_sap3/sap_3_inst.alu_inst.tmp[4] ));
 sg13g2_a22oi_1 \heichips25_sap3/_2880_  (.Y(\heichips25_sap3/_0521_ ),
    .B1(\heichips25_sap3/_0445_ ),
    .B2(\heichips25_sap3/_0356_ ),
    .A2(\heichips25_sap3/_0406_ ),
    .A1(\heichips25_sap3/net154 ));
 sg13g2_xnor2_1 \heichips25_sap3/_2881_  (.Y(\heichips25_sap3/_0522_ ),
    .A(\heichips25_sap3/_0356_ ),
    .B(\heichips25_sap3/_0367_ ));
 sg13g2_xor2_1 \heichips25_sap3/_2882_  (.B(\heichips25_sap3/_0522_ ),
    .A(\heichips25_sap3/_0379_ ),
    .X(\heichips25_sap3/_0523_ ));
 sg13g2_xor2_1 \heichips25_sap3/_2883_  (.B(\heichips25_sap3/_0406_ ),
    .A(\heichips25_sap3/_0405_ ),
    .X(\heichips25_sap3/_0524_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2884_  (.Y(\heichips25_sap3/_0525_ ),
    .B1(\heichips25_sap3/_0417_ ),
    .B2(\heichips25_sap3/net282 ),
    .A2(\heichips25_sap3/_0416_ ),
    .A1(\heichips25_sap3/net278 ));
 sg13g2_o21ai_1 \heichips25_sap3/_2885_  (.B1(\heichips25_sap3/_0525_ ),
    .Y(\heichips25_sap3/_0526_ ),
    .A1(\heichips25_sap3/net280 ),
    .A2(\heichips25_sap3/_0441_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_2886_  (.B2(\heichips25_sap3/_0340_ ),
    .C1(\heichips25_sap3/_0526_ ),
    .B1(\heichips25_sap3/_0524_ ),
    .A1(\heichips25_sap3/_0338_ ),
    .Y(\heichips25_sap3/_0527_ ),
    .A2(\heichips25_sap3/_0523_ ));
 sg13g2_nand4_1 \heichips25_sap3/_2887_  (.B(\heichips25_sap3/_0520_ ),
    .C(\heichips25_sap3/_0521_ ),
    .A(\heichips25_sap3/_0519_ ),
    .Y(\heichips25_sap3/_0528_ ),
    .D(\heichips25_sap3/_0527_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2888_  (.A(\heichips25_sap3/net64 ),
    .B(\heichips25_sap3/_0528_ ),
    .Y(\heichips25_sap3/_0529_ ));
 sg13g2_xnor2_1 \heichips25_sap3/_2889_  (.Y(\heichips25_sap3/_0530_ ),
    .A(\heichips25_sap3/net281 ),
    .B(\heichips25_sap3/net211 ));
 sg13g2_o21ai_1 \heichips25_sap3/_2890_  (.B1(\heichips25_sap3/_0504_ ),
    .Y(\heichips25_sap3/_0531_ ),
    .A1(\heichips25_sap3/_0501_ ),
    .A2(\heichips25_sap3/_0503_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2891_  (.A(\heichips25_sap3/_0530_ ),
    .B(\heichips25_sap3/_0531_ ),
    .Y(\heichips25_sap3/_0532_ ));
 sg13g2_a21o_1 \heichips25_sap3/_2892_  (.A2(\heichips25_sap3/_0531_ ),
    .A1(\heichips25_sap3/_0530_ ),
    .B1(\heichips25_sap3/_1869_ ),
    .X(\heichips25_sap3/_0533_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2893_  (.B1(\heichips25_sap3/_0529_ ),
    .Y(\heichips25_sap3/_0534_ ),
    .A1(\heichips25_sap3/_0532_ ),
    .A2(\heichips25_sap3/_0533_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2894_  (.A1(\heichips25_sap3/net65 ),
    .A2(\heichips25_sap3/_0522_ ),
    .Y(\heichips25_sap3/_0535_ ),
    .B1(\heichips25_sap3/net203 ));
 sg13g2_a221oi_1 \heichips25_sap3/_2895_  (.B2(\heichips25_sap3/_0535_ ),
    .C1(\heichips25_sap3/net157 ),
    .B1(\heichips25_sap3/_0534_ ),
    .A1(\heichips25_sap3/sap_3_inst.alu_inst.act[4] ),
    .Y(\heichips25_sap3/_0536_ ),
    .A2(\heichips25_sap3/net203 ));
 sg13g2_nor3_1 \heichips25_sap3/_2896_  (.A(\heichips25_sap3/net69 ),
    .B(\heichips25_sap3/_0518_ ),
    .C(\heichips25_sap3/_0536_ ),
    .Y(\heichips25_sap3/_0537_ ));
 sg13g2_a21o_1 \heichips25_sap3/_2897_  (.A2(\heichips25_sap3/net69 ),
    .A1(\heichips25_sap3/net281 ),
    .B1(\heichips25_sap3/_0537_ ),
    .X(\heichips25_sap3/_0044_ ));
 sg13g2_nor2b_1 \heichips25_sap3/_2898_  (.A(\uio_out_sap3[5] ),
    .B_N(\heichips25_sap3/net157 ),
    .Y(\heichips25_sap3/_0538_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_2899_  (.Y(\heichips25_sap3/_0539_ ),
    .B(\heichips25_sap3/net159 ),
    .A_N(\heichips25_sap3/_0353_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2900_  (.Y(\heichips25_sap3/_0540_ ),
    .B1(\heichips25_sap3/_0449_ ),
    .B2(\heichips25_sap3/_0351_ ),
    .A2(\heichips25_sap3/_0445_ ),
    .A1(\heichips25_sap3/_0380_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_2901_  (.Y(\heichips25_sap3/_0541_ ),
    .B(\heichips25_sap3/net154 ),
    .A_N(\heichips25_sap3/_0408_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2902_  (.A(\heichips25_sap3/net278 ),
    .B(\heichips25_sap3/_0441_ ),
    .Y(\heichips25_sap3/_0542_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_2903_  (.B2(\heichips25_sap3/net280 ),
    .C1(\heichips25_sap3/_0542_ ),
    .B1(\heichips25_sap3/_0417_ ),
    .A1(\heichips25_sap3/net276 ),
    .Y(\heichips25_sap3/_0543_ ),
    .A2(\heichips25_sap3/_0416_ ));
 sg13g2_nand4_1 \heichips25_sap3/_2904_  (.B(\heichips25_sap3/_0540_ ),
    .C(\heichips25_sap3/_0541_ ),
    .A(\heichips25_sap3/_0539_ ),
    .Y(\heichips25_sap3/_0544_ ),
    .D(\heichips25_sap3/_0543_ ));
 sg13g2_xor2_1 \heichips25_sap3/_2905_  (.B(\heichips25_sap3/_0380_ ),
    .A(\heichips25_sap3/_0368_ ),
    .X(\heichips25_sap3/_0545_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2906_  (.B1(\heichips25_sap3/_0545_ ),
    .Y(\heichips25_sap3/_0546_ ),
    .A1(\heichips25_sap3/_0379_ ),
    .A2(\heichips25_sap3/_0522_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2907_  (.A(\heichips25_sap3/_0379_ ),
    .B(\heichips25_sap3/_0522_ ),
    .C(\heichips25_sap3/_0545_ ),
    .Y(\heichips25_sap3/_0547_ ));
 sg13g2_nand3b_1 \heichips25_sap3/_2908_  (.B(\heichips25_sap3/_0338_ ),
    .C(\heichips25_sap3/_0546_ ),
    .Y(\heichips25_sap3/_0548_ ),
    .A_N(\heichips25_sap3/_0547_ ));
 sg13g2_xor2_1 \heichips25_sap3/_2909_  (.B(\heichips25_sap3/_0408_ ),
    .A(\heichips25_sap3/_0407_ ),
    .X(\heichips25_sap3/_0549_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2910_  (.B1(\heichips25_sap3/_0548_ ),
    .Y(\heichips25_sap3/_0550_ ),
    .A1(\heichips25_sap3/_0341_ ),
    .A2(\heichips25_sap3/_0549_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2911_  (.A(\heichips25_sap3/net65 ),
    .B(\heichips25_sap3/_0544_ ),
    .C(\heichips25_sap3/_0550_ ),
    .Y(\heichips25_sap3/_0551_ ));
 sg13g2_a21o_1 \heichips25_sap3/_2912_  (.A2(\heichips25_sap3/net211 ),
    .A1(\heichips25_sap3/net281 ),
    .B1(\heichips25_sap3/_0532_ ),
    .X(\heichips25_sap3/_0552_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2913_  (.Y(\heichips25_sap3/_0553_ ),
    .A(\heichips25_sap3/net278 ),
    .B(\heichips25_sap3/net211 ));
 sg13g2_xnor2_1 \heichips25_sap3/_2914_  (.Y(\heichips25_sap3/_0554_ ),
    .A(\heichips25_sap3/_1382_ ),
    .B(\heichips25_sap3/net211 ));
 sg13g2_xnor2_1 \heichips25_sap3/_2915_  (.Y(\heichips25_sap3/_0555_ ),
    .A(\heichips25_sap3/_0552_ ),
    .B(\heichips25_sap3/_0554_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2916_  (.B1(\heichips25_sap3/_0551_ ),
    .Y(\heichips25_sap3/_0556_ ),
    .A1(\heichips25_sap3/_1869_ ),
    .A2(\heichips25_sap3/_0555_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2917_  (.A1(\heichips25_sap3/net65 ),
    .A2(\heichips25_sap3/_0545_ ),
    .Y(\heichips25_sap3/_0557_ ),
    .B1(\heichips25_sap3/net203 ));
 sg13g2_a221oi_1 \heichips25_sap3/_2918_  (.B2(\heichips25_sap3/_0557_ ),
    .C1(\heichips25_sap3/net157 ),
    .B1(\heichips25_sap3/_0556_ ),
    .A1(\heichips25_sap3/sap_3_inst.alu_inst.act[5] ),
    .Y(\heichips25_sap3/_0558_ ),
    .A2(\heichips25_sap3/net203 ));
 sg13g2_nor3_1 \heichips25_sap3/_2919_  (.A(\heichips25_sap3/net69 ),
    .B(\heichips25_sap3/_0538_ ),
    .C(\heichips25_sap3/_0558_ ),
    .Y(\heichips25_sap3/_0559_ ));
 sg13g2_a21o_1 \heichips25_sap3/_2920_  (.A2(\heichips25_sap3/net69 ),
    .A1(\heichips25_sap3/net279 ),
    .B1(\heichips25_sap3/_0559_ ),
    .X(\heichips25_sap3/_0045_ ));
 sg13g2_nor2b_1 \heichips25_sap3/_2921_  (.A(net43),
    .B_N(\heichips25_sap3/net157 ),
    .Y(\heichips25_sap3/_0560_ ));
 sg13g2_xor2_1 \heichips25_sap3/_2922_  (.B(\heichips25_sap3/_0369_ ),
    .A(\heichips25_sap3/_0350_ ),
    .X(\heichips25_sap3/_0561_ ));
 sg13g2_inv_1 \heichips25_sap3/_2923_  (.Y(\heichips25_sap3/_0562_ ),
    .A(\heichips25_sap3/_0561_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2924_  (.Y(\heichips25_sap3/_0563_ ),
    .A(\heichips25_sap3/_0547_ ),
    .B(\heichips25_sap3/_0561_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2925_  (.B1(\heichips25_sap3/_0338_ ),
    .Y(\heichips25_sap3/_0564_ ),
    .A1(\heichips25_sap3/_0547_ ),
    .A2(\heichips25_sap3/_0561_ ));
 sg13g2_nor2b_1 \heichips25_sap3/_2926_  (.A(\heichips25_sap3/_0564_ ),
    .B_N(\heichips25_sap3/_0563_ ),
    .Y(\heichips25_sap3/_0565_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2927_  (.Y(\heichips25_sap3/_0566_ ),
    .A(\heichips25_sap3/net278 ),
    .B(\heichips25_sap3/_0417_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2928_  (.Y(\heichips25_sap3/_0567_ ),
    .B1(\heichips25_sap3/_0449_ ),
    .B2(\heichips25_sap3/_0349_ ),
    .A2(\heichips25_sap3/_0416_ ),
    .A1(\heichips25_sap3/net274 ));
 sg13g2_nand2_1 \heichips25_sap3/_2929_  (.Y(\heichips25_sap3/_0568_ ),
    .A(\heichips25_sap3/_0350_ ),
    .B(\heichips25_sap3/_0445_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2930_  (.B1(\heichips25_sap3/net159 ),
    .Y(\heichips25_sap3/_0569_ ),
    .A1(\heichips25_sap3/net276 ),
    .A2(\heichips25_sap3/sap_3_inst.alu_inst.tmp[6] ));
 sg13g2_nand4_1 \heichips25_sap3/_2931_  (.B(\heichips25_sap3/_0567_ ),
    .C(\heichips25_sap3/_0568_ ),
    .A(\heichips25_sap3/_0566_ ),
    .Y(\heichips25_sap3/_0570_ ),
    .D(\heichips25_sap3/_0569_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_2932_  (.B2(\heichips25_sap3/_1384_ ),
    .C1(\heichips25_sap3/_0570_ ),
    .B1(\heichips25_sap3/_0442_ ),
    .A1(\heichips25_sap3/_0343_ ),
    .Y(\heichips25_sap3/_0571_ ),
    .A2(\heichips25_sap3/_0399_ ));
 sg13g2_xor2_1 \heichips25_sap3/_2933_  (.B(\heichips25_sap3/_0409_ ),
    .A(\heichips25_sap3/_0399_ ),
    .X(\heichips25_sap3/_0572_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2934_  (.B1(\heichips25_sap3/_0571_ ),
    .Y(\heichips25_sap3/_0573_ ),
    .A1(\heichips25_sap3/_0341_ ),
    .A2(\heichips25_sap3/_0572_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2935_  (.A(\heichips25_sap3/net65 ),
    .B(\heichips25_sap3/_0565_ ),
    .C(\heichips25_sap3/_0573_ ),
    .Y(\heichips25_sap3/_0574_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2936_  (.Y(\heichips25_sap3/_0575_ ),
    .A(\heichips25_sap3/net276 ),
    .B(\heichips25_sap3/net211 ));
 sg13g2_xnor2_1 \heichips25_sap3/_2937_  (.Y(\heichips25_sap3/_0576_ ),
    .A(\heichips25_sap3/net276 ),
    .B(\heichips25_sap3/net211 ));
 sg13g2_o21ai_1 \heichips25_sap3/_2938_  (.B1(\heichips25_sap3/_0552_ ),
    .Y(\heichips25_sap3/_0577_ ),
    .A1(\heichips25_sap3/net279 ),
    .A2(\heichips25_sap3/net211 ));
 sg13g2_and2_1 \heichips25_sap3/_2939_  (.A(\heichips25_sap3/_0553_ ),
    .B(\heichips25_sap3/_0577_ ),
    .X(\heichips25_sap3/_0578_ ));
 sg13g2_xnor2_1 \heichips25_sap3/_2940_  (.Y(\heichips25_sap3/_0579_ ),
    .A(\heichips25_sap3/_0576_ ),
    .B(\heichips25_sap3/_0578_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2941_  (.B1(\heichips25_sap3/_0574_ ),
    .Y(\heichips25_sap3/_0580_ ),
    .A1(\heichips25_sap3/_1869_ ),
    .A2(\heichips25_sap3/_0579_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2942_  (.A1(\heichips25_sap3/net65 ),
    .A2(\heichips25_sap3/_0562_ ),
    .Y(\heichips25_sap3/_0581_ ),
    .B1(\heichips25_sap3/net203 ));
 sg13g2_a221oi_1 \heichips25_sap3/_2943_  (.B2(\heichips25_sap3/_0581_ ),
    .C1(\heichips25_sap3/net157 ),
    .B1(\heichips25_sap3/_0580_ ),
    .A1(\heichips25_sap3/sap_3_inst.alu_inst.act[6] ),
    .Y(\heichips25_sap3/_0582_ ),
    .A2(\heichips25_sap3/net203 ));
 sg13g2_nor3_1 \heichips25_sap3/_2944_  (.A(\heichips25_sap3/net69 ),
    .B(\heichips25_sap3/_0560_ ),
    .C(\heichips25_sap3/_0582_ ),
    .Y(\heichips25_sap3/_0583_ ));
 sg13g2_a21o_1 \heichips25_sap3/_2945_  (.A2(\heichips25_sap3/net69 ),
    .A1(\heichips25_sap3/net277 ),
    .B1(\heichips25_sap3/_0583_ ),
    .X(\heichips25_sap3/_0046_ ));
 sg13g2_nor2b_1 \heichips25_sap3/_2946_  (.A(net47),
    .B_N(\heichips25_sap3/_0434_ ),
    .Y(\heichips25_sap3/_0584_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2947_  (.B1(\heichips25_sap3/_0575_ ),
    .Y(\heichips25_sap3/_0585_ ),
    .A1(\heichips25_sap3/_0576_ ),
    .A2(\heichips25_sap3/_0578_ ));
 sg13g2_xnor2_1 \heichips25_sap3/_2948_  (.Y(\heichips25_sap3/_0586_ ),
    .A(\heichips25_sap3/_1374_ ),
    .B(\heichips25_sap3/net212 ));
 sg13g2_xnor2_1 \heichips25_sap3/_2949_  (.Y(\heichips25_sap3/_0587_ ),
    .A(\heichips25_sap3/_0585_ ),
    .B(\heichips25_sap3/_0586_ ));
 sg13g2_xor2_1 \heichips25_sap3/_2950_  (.B(\heichips25_sap3/_0381_ ),
    .A(\heichips25_sap3/_0370_ ),
    .X(\heichips25_sap3/_0588_ ));
 sg13g2_xor2_1 \heichips25_sap3/_2951_  (.B(\heichips25_sap3/_0588_ ),
    .A(\heichips25_sap3/_0563_ ),
    .X(\heichips25_sap3/_0589_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_2952_  (.Y(\heichips25_sap3/_0590_ ),
    .B(\heichips25_sap3/_0449_ ),
    .A_N(\heichips25_sap3/_0348_ ));
 sg13g2_nand3_1 \heichips25_sap3/_2953_  (.B(\heichips25_sap3/_1892_ ),
    .C(\heichips25_sap3/_1896_ ),
    .A(\heichips25_sap3/net254 ),
    .Y(\heichips25_sap3/_0591_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2954_  (.Y(\heichips25_sap3/_0592_ ),
    .A(\heichips25_sap3/_1374_ ),
    .B(\heichips25_sap3/_0442_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_2955_  (.Y(\heichips25_sap3/_0593_ ),
    .B(\heichips25_sap3/_1895_ ),
    .A_N(\heichips25_sap3/_0347_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2956_  (.Y(\heichips25_sap3/_0594_ ),
    .A(\heichips25_sap3/_0590_ ),
    .B(\heichips25_sap3/_0593_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_2957_  (.B2(\heichips25_sap3/_0381_ ),
    .C1(\heichips25_sap3/_0594_ ),
    .B1(\heichips25_sap3/_0445_ ),
    .A1(\heichips25_sap3/net276 ),
    .Y(\heichips25_sap3/_0595_ ),
    .A2(\heichips25_sap3/_0417_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2958_  (.A1(\heichips25_sap3/_0343_ ),
    .A2(\heichips25_sap3/_0412_ ),
    .Y(\heichips25_sap3/_0596_ ),
    .B1(\heichips25_sap3/net65 ));
 sg13g2_nand4_1 \heichips25_sap3/_2959_  (.B(\heichips25_sap3/_0592_ ),
    .C(\heichips25_sap3/_0595_ ),
    .A(\heichips25_sap3/_0591_ ),
    .Y(\heichips25_sap3/_0597_ ),
    .D(\heichips25_sap3/_0596_ ));
 sg13g2_xor2_1 \heichips25_sap3/_2960_  (.B(\heichips25_sap3/_0412_ ),
    .A(\heichips25_sap3/_0410_ ),
    .X(\heichips25_sap3/_0598_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_2961_  (.B2(\heichips25_sap3/_0340_ ),
    .C1(\heichips25_sap3/_0597_ ),
    .B1(\heichips25_sap3/_0598_ ),
    .A1(\heichips25_sap3/_0338_ ),
    .Y(\heichips25_sap3/_0599_ ),
    .A2(\heichips25_sap3/_0589_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2962_  (.B1(\heichips25_sap3/_0599_ ),
    .Y(\heichips25_sap3/_0600_ ),
    .A1(\heichips25_sap3/_1869_ ),
    .A2(\heichips25_sap3/_0587_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2963_  (.A1(\heichips25_sap3/net65 ),
    .A2(\heichips25_sap3/_0588_ ),
    .Y(\heichips25_sap3/_0601_ ),
    .B1(\heichips25_sap3/_0436_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_2964_  (.B2(\heichips25_sap3/_0601_ ),
    .C1(\heichips25_sap3/_0434_ ),
    .B1(\heichips25_sap3/_0600_ ),
    .A1(\heichips25_sap3/sap_3_inst.alu_inst.act[7] ),
    .Y(\heichips25_sap3/_0602_ ),
    .A2(\heichips25_sap3/_0436_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2965_  (.A(\heichips25_sap3/_0440_ ),
    .B(\heichips25_sap3/_0584_ ),
    .C(\heichips25_sap3/_0602_ ),
    .Y(\heichips25_sap3/_0603_ ));
 sg13g2_a21o_1 \heichips25_sap3/_2966_  (.A2(\heichips25_sap3/net70 ),
    .A1(\heichips25_sap3/net275 ),
    .B1(\heichips25_sap3/_0603_ ),
    .X(\heichips25_sap3/_0047_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2967_  (.Y(\heichips25_sap3/_0604_ ),
    .A(\heichips25_sap3/_1641_ ),
    .B(\heichips25_sap3/_1646_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_2968_  (.B1(\heichips25_sap3/_1767_ ),
    .Y(\heichips25_sap3/_0605_ ),
    .A1(\heichips25_sap3/_0426_ ),
    .A2(\heichips25_sap3/_0604_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2969_  (.A(\heichips25_sap3/_1883_ ),
    .B(\heichips25_sap3/_1893_ ),
    .Y(\heichips25_sap3/_0606_ ));
 sg13g2_nor2_1 \heichips25_sap3/_2970_  (.A(\heichips25_sap3/net167 ),
    .B(\heichips25_sap3/net153 ),
    .Y(\heichips25_sap3/_0607_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2971_  (.Y(\heichips25_sap3/_0608_ ),
    .A(\heichips25_sap3/sap_3_inst.alu_inst.act[0] ),
    .B(\heichips25_sap3/_0607_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2972_  (.Y(\heichips25_sap3/_0609_ ),
    .B1(\heichips25_sap3/net153 ),
    .B2(\heichips25_sap3/_0372_ ),
    .A2(\heichips25_sap3/net167 ),
    .A1(\heichips25_sap3/sap_3_inst.alu_inst.acc[0] ));
 sg13g2_nand2_1 \heichips25_sap3/_2973_  (.Y(\heichips25_sap3/_0048_ ),
    .A(\heichips25_sap3/_0608_ ),
    .B(\heichips25_sap3/_0609_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2974_  (.Y(\heichips25_sap3/_0610_ ),
    .A(\heichips25_sap3/sap_3_inst.alu_inst.act[1] ),
    .B(\heichips25_sap3/_0607_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2975_  (.Y(\heichips25_sap3/_0611_ ),
    .B1(\heichips25_sap3/net153 ),
    .B2(\heichips25_sap3/_0400_ ),
    .A2(\heichips25_sap3/net167 ),
    .A1(\heichips25_sap3/net286 ));
 sg13g2_nand2_1 \heichips25_sap3/_2976_  (.Y(\heichips25_sap3/_0049_ ),
    .A(\heichips25_sap3/_0610_ ),
    .B(\heichips25_sap3/_0611_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2977_  (.Y(\heichips25_sap3/_0612_ ),
    .A(\heichips25_sap3/sap_3_inst.alu_inst.act[2] ),
    .B(\heichips25_sap3/_0607_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2978_  (.Y(\heichips25_sap3/_0613_ ),
    .B1(\heichips25_sap3/net153 ),
    .B2(\heichips25_sap3/_0403_ ),
    .A2(\heichips25_sap3/net167 ),
    .A1(\heichips25_sap3/net284 ));
 sg13g2_nand2_1 \heichips25_sap3/_2979_  (.Y(\heichips25_sap3/_0050_ ),
    .A(\heichips25_sap3/_0612_ ),
    .B(\heichips25_sap3/_0613_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2980_  (.Y(\heichips25_sap3/_0614_ ),
    .A(\heichips25_sap3/sap_3_inst.alu_inst.act[3] ),
    .B(\heichips25_sap3/_0607_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2981_  (.Y(\heichips25_sap3/_0615_ ),
    .B1(\heichips25_sap3/net153 ),
    .B2(\heichips25_sap3/_0404_ ),
    .A2(\heichips25_sap3/net167 ),
    .A1(\heichips25_sap3/net282 ));
 sg13g2_nand2_1 \heichips25_sap3/_2982_  (.Y(\heichips25_sap3/_0051_ ),
    .A(\heichips25_sap3/_0614_ ),
    .B(\heichips25_sap3/_0615_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2983_  (.Y(\heichips25_sap3/_0616_ ),
    .A(\heichips25_sap3/sap_3_inst.alu_inst.act[4] ),
    .B(\heichips25_sap3/_0607_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2984_  (.Y(\heichips25_sap3/_0617_ ),
    .B1(\heichips25_sap3/net153 ),
    .B2(\heichips25_sap3/_0406_ ),
    .A2(\heichips25_sap3/net167 ),
    .A1(\heichips25_sap3/net281 ));
 sg13g2_nand2_1 \heichips25_sap3/_2985_  (.Y(\heichips25_sap3/_0052_ ),
    .A(\heichips25_sap3/_0616_ ),
    .B(\heichips25_sap3/_0617_ ));
 sg13g2_nor3_1 \heichips25_sap3/_2986_  (.A(\heichips25_sap3/sap_3_inst.alu_inst.act[5] ),
    .B(\heichips25_sap3/net167 ),
    .C(\heichips25_sap3/net153 ),
    .Y(\heichips25_sap3/_0618_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_2987_  (.B2(\heichips25_sap3/_0408_ ),
    .C1(\heichips25_sap3/_0618_ ),
    .B1(\heichips25_sap3/net153 ),
    .A1(\heichips25_sap3/_1382_ ),
    .Y(\heichips25_sap3/_0053_ ),
    .A2(\heichips25_sap3/net167 ));
 sg13g2_nand2_1 \heichips25_sap3/_2988_  (.Y(\heichips25_sap3/_0619_ ),
    .A(\heichips25_sap3/net277 ),
    .B(\heichips25_sap3/_0605_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2989_  (.Y(\heichips25_sap3/_0620_ ),
    .B1(\heichips25_sap3/_0607_ ),
    .B2(\heichips25_sap3/sap_3_inst.alu_inst.act[6] ),
    .A2(\heichips25_sap3/_0606_ ),
    .A1(\heichips25_sap3/_0399_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2990_  (.Y(\heichips25_sap3/_0054_ ),
    .A(\heichips25_sap3/_0619_ ),
    .B(\heichips25_sap3/_0620_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2991_  (.Y(\heichips25_sap3/_0621_ ),
    .A(\heichips25_sap3/sap_3_inst.alu_inst.act[7] ),
    .B(\heichips25_sap3/_0607_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2992_  (.Y(\heichips25_sap3/_0622_ ),
    .B1(\heichips25_sap3/_0606_ ),
    .B2(\heichips25_sap3/_0412_ ),
    .A2(\heichips25_sap3/_0605_ ),
    .A1(\heichips25_sap3/net275 ));
 sg13g2_nand2_1 \heichips25_sap3/_2993_  (.Y(\heichips25_sap3/_0055_ ),
    .A(\heichips25_sap3/_0621_ ),
    .B(\heichips25_sap3/_0622_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2994_  (.A1(\heichips25_sap3/net238 ),
    .A2(\heichips25_sap3/_1614_ ),
    .Y(\heichips25_sap3/_0623_ ),
    .B1(\heichips25_sap3/_1662_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_2995_  (.Y(\heichips25_sap3/_0624_ ),
    .B1(\heichips25_sap3/_1760_ ),
    .B2(\heichips25_sap3/_0623_ ),
    .A2(\heichips25_sap3/_1709_ ),
    .A1(\heichips25_sap3/net224 ));
 sg13g2_nor2_1 \heichips25_sap3/_2996_  (.A(\heichips25_sap3/sap_3_inst.alu_inst.tmp[0] ),
    .B(\heichips25_sap3/net201 ),
    .Y(\heichips25_sap3/_0625_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_2997_  (.A1(\heichips25_sap3/_0212_ ),
    .A2(\heichips25_sap3/net201 ),
    .Y(\heichips25_sap3/_0056_ ),
    .B1(\heichips25_sap3/_0625_ ));
 sg13g2_nand2_1 \heichips25_sap3/_2998_  (.Y(\heichips25_sap3/_0626_ ),
    .A(\uio_out_sap3[1] ),
    .B(\heichips25_sap3/net201 ));
 sg13g2_o21ai_1 \heichips25_sap3/_2999_  (.B1(\heichips25_sap3/_0626_ ),
    .Y(\heichips25_sap3/_0057_ ),
    .A1(\heichips25_sap3/_1396_ ),
    .A2(\heichips25_sap3/net201 ));
 sg13g2_nand2_1 \heichips25_sap3/_3000_  (.Y(\heichips25_sap3/_0627_ ),
    .A(net44),
    .B(\heichips25_sap3/net201 ));
 sg13g2_o21ai_1 \heichips25_sap3/_3001_  (.B1(\heichips25_sap3/_0627_ ),
    .Y(\heichips25_sap3/_0058_ ),
    .A1(\heichips25_sap3/_1397_ ),
    .A2(\heichips25_sap3/net201 ));
 sg13g2_nor2_1 \heichips25_sap3/_3002_  (.A(\heichips25_sap3/sap_3_inst.alu_inst.tmp[3] ),
    .B(\heichips25_sap3/net201 ),
    .Y(\heichips25_sap3/_0628_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3003_  (.A1(\heichips25_sap3/net45 ),
    .A2(\heichips25_sap3/net201 ),
    .Y(\heichips25_sap3/_0059_ ),
    .B1(\heichips25_sap3/_0628_ ));
 sg13g2_mux2_1 \heichips25_sap3/_3004_  (.A0(\heichips25_sap3/sap_3_inst.alu_inst.tmp[4] ),
    .A1(net46),
    .S(\heichips25_sap3/net202 ),
    .X(\heichips25_sap3/_0060_ ));
 sg13g2_mux2_1 \heichips25_sap3/_3005_  (.A0(\heichips25_sap3/sap_3_inst.alu_inst.tmp[5] ),
    .A1(\uio_out_sap3[5] ),
    .S(\heichips25_sap3/net202 ),
    .X(\heichips25_sap3/_0061_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3006_  (.Y(\heichips25_sap3/_0629_ ),
    .A(\heichips25_sap3/net826 ),
    .B(\heichips25_sap3/net202 ));
 sg13g2_o21ai_1 \heichips25_sap3/_3007_  (.B1(\heichips25_sap3/_0629_ ),
    .Y(\heichips25_sap3/_0062_ ),
    .A1(\heichips25_sap3/_1398_ ),
    .A2(\heichips25_sap3/net202 ));
 sg13g2_nand2_1 \heichips25_sap3/_3008_  (.Y(\heichips25_sap3/_0630_ ),
    .A(net47),
    .B(\heichips25_sap3/net202 ));
 sg13g2_o21ai_1 \heichips25_sap3/_3009_  (.B1(\heichips25_sap3/_0630_ ),
    .Y(\heichips25_sap3/_0063_ ),
    .A1(\heichips25_sap3/_1399_ ),
    .A2(\heichips25_sap3/net202 ));
 sg13g2_nand2_1 \heichips25_sap3/_3010_  (.Y(\heichips25_sap3/_0631_ ),
    .A(\heichips25_sap3/net273 ),
    .B(\heichips25_sap3/net231 ));
 sg13g2_o21ai_1 \heichips25_sap3/_3011_  (.B1(\heichips25_sap3/_0631_ ),
    .Y(\heichips25_sap3/_0064_ ),
    .A1(\heichips25_sap3/net231 ),
    .A2(\heichips25_sap3/_0212_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3012_  (.Y(\heichips25_sap3/_0632_ ),
    .A(\heichips25_sap3/net270 ),
    .B(\heichips25_sap3/net231 ));
 sg13g2_o21ai_1 \heichips25_sap3/_3013_  (.B1(\heichips25_sap3/_0632_ ),
    .Y(\heichips25_sap3/_0065_ ),
    .A1(\heichips25_sap3/net233 ),
    .A2(\heichips25_sap3/_1922_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3014_  (.A(\heichips25_sap3/net233 ),
    .B(\uio_out_sap3[2] ),
    .Y(\heichips25_sap3/_0633_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3015_  (.A1(\heichips25_sap3/_1362_ ),
    .A2(\heichips25_sap3/net231 ),
    .Y(\heichips25_sap3/_0066_ ),
    .B1(\heichips25_sap3/_0633_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3016_  (.Y(\heichips25_sap3/_0634_ ),
    .A(\heichips25_sap3/net265 ),
    .B(\heichips25_sap3/net232 ));
 sg13g2_o21ai_1 \heichips25_sap3/_3017_  (.B1(\heichips25_sap3/_0634_ ),
    .Y(\heichips25_sap3/_0067_ ),
    .A1(\heichips25_sap3/net232 ),
    .A2(\heichips25_sap3/_0242_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3018_  (.A(\heichips25_sap3/net232 ),
    .B(\uio_out_sap3[4] ),
    .Y(\heichips25_sap3/_0635_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3019_  (.A1(\heichips25_sap3/_1364_ ),
    .A2(\heichips25_sap3/net232 ),
    .Y(\heichips25_sap3/_0068_ ),
    .B1(\heichips25_sap3/_0635_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3020_  (.A(\heichips25_sap3/net233 ),
    .B(\uio_out_sap3[5] ),
    .Y(\heichips25_sap3/_0636_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3021_  (.A1(\heichips25_sap3/_1365_ ),
    .A2(\heichips25_sap3/net233 ),
    .Y(\heichips25_sap3/_0069_ ),
    .B1(\heichips25_sap3/_0636_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3022_  (.A(\heichips25_sap3/net231 ),
    .B(\heichips25_sap3/net826 ),
    .Y(\heichips25_sap3/_0637_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3023_  (.A1(\heichips25_sap3/_1361_ ),
    .A2(\heichips25_sap3/net231 ),
    .Y(\heichips25_sap3/_0070_ ),
    .B1(\heichips25_sap3/_0637_ ));
 sg13g2_mux2_1 \heichips25_sap3/_3024_  (.A0(\uio_out_sap3[7] ),
    .A1(\heichips25_sap3/net259 ),
    .S(\heichips25_sap3/net231 ),
    .X(\heichips25_sap3/_0071_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3025_  (.A1(\heichips25_sap3/net235 ),
    .A2(\heichips25_sap3/net229 ),
    .Y(\heichips25_sap3/_0638_ ),
    .B1(\heichips25_sap3/_1492_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_3026_  (.B2(\heichips25_sap3/_1541_ ),
    .C1(\heichips25_sap3/_0638_ ),
    .B1(\heichips25_sap3/_1759_ ),
    .A1(\heichips25_sap3/_1494_ ),
    .Y(\heichips25_sap3/_0639_ ),
    .A2(\heichips25_sap3/_1626_ ));
 sg13g2_nor3_1 \heichips25_sap3/_3027_  (.A(\heichips25_sap3/_1525_ ),
    .B(\heichips25_sap3/_1535_ ),
    .C(\heichips25_sap3/_0639_ ),
    .Y(\heichips25_sap3/_0640_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3028_  (.A(\heichips25_sap3/_1520_ ),
    .B(\heichips25_sap3/_1658_ ),
    .Y(\heichips25_sap3/_0641_ ));
 sg13g2_nand4_1 \heichips25_sap3/_3029_  (.B(\heichips25_sap3/_1521_ ),
    .C(\heichips25_sap3/_1527_ ),
    .A(\heichips25_sap3/_1504_ ),
    .Y(\heichips25_sap3/_0642_ ),
    .D(\heichips25_sap3/_1565_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3030_  (.A1(\heichips25_sap3/_1485_ ),
    .A2(\heichips25_sap3/_0642_ ),
    .Y(\heichips25_sap3/_0643_ ),
    .B1(\heichips25_sap3/_1697_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3031_  (.A(\heichips25_sap3/_1527_ ),
    .B(\heichips25_sap3/_1569_ ),
    .Y(\heichips25_sap3/_0644_ ));
 sg13g2_nor3_1 \heichips25_sap3/_3032_  (.A(\heichips25_sap3/_1475_ ),
    .B(\heichips25_sap3/net226 ),
    .C(\heichips25_sap3/_1643_ ),
    .Y(\heichips25_sap3/_0645_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3033_  (.Y(\heichips25_sap3/_0646_ ),
    .A(\heichips25_sap3/_1644_ ),
    .B(\heichips25_sap3/_1762_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3034_  (.B1(\heichips25_sap3/net263 ),
    .Y(\heichips25_sap3/_0647_ ),
    .A1(\heichips25_sap3/_0644_ ),
    .A2(\heichips25_sap3/_0645_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3035_  (.A1(\heichips25_sap3/_1486_ ),
    .A2(\heichips25_sap3/_1572_ ),
    .Y(\heichips25_sap3/_0648_ ),
    .B1(\heichips25_sap3/_1510_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3036_  (.Y(\heichips25_sap3/_0649_ ),
    .B1(\heichips25_sap3/_1580_ ),
    .B2(\heichips25_sap3/_1486_ ),
    .A2(\heichips25_sap3/_1532_ ),
    .A1(\heichips25_sap3/_1513_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3037_  (.Y(\heichips25_sap3/_0650_ ),
    .A(\heichips25_sap3/_1486_ ),
    .B(\heichips25_sap3/_1625_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_3038_  (.B2(\heichips25_sap3/_1664_ ),
    .C1(\heichips25_sap3/_0648_ ),
    .B1(\heichips25_sap3/_0650_ ),
    .A1(\heichips25_sap3/net263 ),
    .Y(\heichips25_sap3/_0651_ ),
    .A2(\heichips25_sap3/_1773_ ));
 sg13g2_nor3_1 \heichips25_sap3/_3039_  (.A(\heichips25_sap3/net220 ),
    .B(\heichips25_sap3/_1778_ ),
    .C(\heichips25_sap3/_0649_ ),
    .Y(\heichips25_sap3/_0652_ ));
 sg13g2_nand4_1 \heichips25_sap3/_3040_  (.B(\heichips25_sap3/_0647_ ),
    .C(\heichips25_sap3/_0651_ ),
    .A(\heichips25_sap3/_0643_ ),
    .Y(\heichips25_sap3/_0653_ ),
    .D(\heichips25_sap3/_0652_ ));
 sg13g2_nor3_1 \heichips25_sap3/_3041_  (.A(\heichips25_sap3/net234 ),
    .B(\heichips25_sap3/_1501_ ),
    .C(\heichips25_sap3/_1506_ ),
    .Y(\heichips25_sap3/_0654_ ));
 sg13g2_nor3_1 \heichips25_sap3/_3042_  (.A(\heichips25_sap3/_1450_ ),
    .B(\heichips25_sap3/net234 ),
    .C(\heichips25_sap3/_1643_ ),
    .Y(\heichips25_sap3/_0655_ ));
 sg13g2_nand3_1 \heichips25_sap3/_3043_  (.B(\heichips25_sap3/net238 ),
    .C(\heichips25_sap3/_1644_ ),
    .A(\heichips25_sap3/_1449_ ),
    .Y(\heichips25_sap3/_0656_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3044_  (.B1(\heichips25_sap3/net263 ),
    .Y(\heichips25_sap3/_0657_ ),
    .A1(\heichips25_sap3/_0654_ ),
    .A2(\heichips25_sap3/_0655_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3045_  (.A1(\heichips25_sap3/net220 ),
    .A2(\heichips25_sap3/_0657_ ),
    .Y(\heichips25_sap3/_0658_ ),
    .B1(\heichips25_sap3/net248 ));
 sg13g2_o21ai_1 \heichips25_sap3/_3046_  (.B1(\heichips25_sap3/_0658_ ),
    .Y(\heichips25_sap3/_0659_ ),
    .A1(\heichips25_sap3/_0640_ ),
    .A2(\heichips25_sap3/_0653_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3047_  (.Y(\heichips25_sap3/_0660_ ),
    .A(\heichips25_sap3/_1364_ ),
    .B(\heichips25_sap3/_1451_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3048_  (.A1(\heichips25_sap3/net227 ),
    .A2(\heichips25_sap3/_1644_ ),
    .Y(\heichips25_sap3/_0661_ ),
    .B1(\heichips25_sap3/net241 ));
 sg13g2_nor3_1 \heichips25_sap3/_3049_  (.A(\heichips25_sap3/_1455_ ),
    .B(\heichips25_sap3/_1465_ ),
    .C(\heichips25_sap3/_0661_ ),
    .Y(\heichips25_sap3/_0662_ ));
 sg13g2_inv_1 \heichips25_sap3/_3050_  (.Y(\heichips25_sap3/_0663_ ),
    .A(\heichips25_sap3/_0662_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3051_  (.Y(\heichips25_sap3/_0664_ ),
    .A(\heichips25_sap3/_0660_ ),
    .B(\heichips25_sap3/_0662_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3052_  (.A1(\heichips25_sap3/net241 ),
    .A2(\heichips25_sap3/_0659_ ),
    .Y(\heichips25_sap3/_0665_ ),
    .B1(\heichips25_sap3/_0663_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3053_  (.A1(\heichips25_sap3/net241 ),
    .A2(\heichips25_sap3/_0659_ ),
    .Y(\heichips25_sap3/_0666_ ),
    .B1(\heichips25_sap3/_0664_ ));
 sg13g2_a21o_1 \heichips25_sap3/_3054_  (.A2(\heichips25_sap3/_0659_ ),
    .A1(\heichips25_sap3/net241 ),
    .B1(\heichips25_sap3/_0664_ ),
    .X(\heichips25_sap3/_0667_ ));
 sg13g2_or2_1 \heichips25_sap3/_3055_  (.X(\heichips25_sap3/_0668_ ),
    .B(\heichips25_sap3/_1725_ ),
    .A(\heichips25_sap3/_1363_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3056_  (.A(\heichips25_sap3/_1441_ ),
    .B(\heichips25_sap3/_1495_ ),
    .Y(\heichips25_sap3/_0669_ ));
 sg13g2_nor4_1 \heichips25_sap3/_3057_  (.A(\heichips25_sap3/net245 ),
    .B(\heichips25_sap3/_1515_ ),
    .C(\heichips25_sap3/_1537_ ),
    .D(\heichips25_sap3/_0669_ ),
    .Y(\heichips25_sap3/_0670_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3058_  (.Y(\heichips25_sap3/_0671_ ),
    .B1(\heichips25_sap3/_0670_ ),
    .B2(\heichips25_sap3/_0641_ ),
    .A2(\heichips25_sap3/_0668_ ),
    .A1(\heichips25_sap3/net225 ));
 sg13g2_nand3_1 \heichips25_sap3/_3059_  (.B(\heichips25_sap3/net239 ),
    .C(\heichips25_sap3/_1721_ ),
    .A(\heichips25_sap3/_1449_ ),
    .Y(\heichips25_sap3/_0672_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3060_  (.Y(\heichips25_sap3/_0673_ ),
    .A(\heichips25_sap3/net266 ),
    .B(\heichips25_sap3/_1773_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3061_  (.Y(\heichips25_sap3/_0674_ ),
    .B1(\heichips25_sap3/_1605_ ),
    .B2(\heichips25_sap3/_1664_ ),
    .A2(\heichips25_sap3/_1517_ ),
    .A1(\heichips25_sap3/_1496_ ));
 sg13g2_nand3_1 \heichips25_sap3/_3062_  (.B(\heichips25_sap3/_0673_ ),
    .C(\heichips25_sap3/_0674_ ),
    .A(\heichips25_sap3/_0672_ ),
    .Y(\heichips25_sap3/_0675_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3063_  (.B1(\heichips25_sap3/net241 ),
    .Y(\heichips25_sap3/_0676_ ),
    .A1(\heichips25_sap3/_0671_ ),
    .A2(\heichips25_sap3/_0675_ ));
 sg13g2_or4_1 \heichips25_sap3/_3064_  (.A(\heichips25_sap3/net258 ),
    .B(\heichips25_sap3/_1448_ ),
    .C(\heichips25_sap3/net226 ),
    .D(\heichips25_sap3/_1722_ ),
    .X(\heichips25_sap3/_0677_ ));
 sg13g2_and2_1 \heichips25_sap3/_3065_  (.A(\heichips25_sap3/_0676_ ),
    .B(\heichips25_sap3/_0677_ ),
    .X(\heichips25_sap3/_0678_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3066_  (.Y(\heichips25_sap3/_0679_ ),
    .A(\heichips25_sap3/_0676_ ),
    .B(\heichips25_sap3/_0677_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3067_  (.A(\heichips25_sap3/_0666_ ),
    .B(\heichips25_sap3/_0679_ ),
    .Y(\heichips25_sap3/_0680_ ));
 sg13g2_nand3_1 \heichips25_sap3/_3068_  (.B(\heichips25_sap3/_1526_ ),
    .C(\heichips25_sap3/_1568_ ),
    .A(\heichips25_sap3/_1507_ ),
    .Y(\heichips25_sap3/_0681_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3069_  (.Y(\heichips25_sap3/_0682_ ),
    .B1(\heichips25_sap3/_0681_ ),
    .B2(\heichips25_sap3/_1486_ ),
    .A2(\heichips25_sap3/_1754_ ),
    .A1(\heichips25_sap3/_1685_ ));
 sg13g2_nor3_1 \heichips25_sap3/_3070_  (.A(\heichips25_sap3/_1365_ ),
    .B(\heichips25_sap3/_1480_ ),
    .C(\heichips25_sap3/_1619_ ),
    .Y(\heichips25_sap3/_0683_ ));
 sg13g2_nand3_1 \heichips25_sap3/_3071_  (.B(\heichips25_sap3/net228 ),
    .C(\heichips25_sap3/_1668_ ),
    .A(\heichips25_sap3/_1474_ ),
    .Y(\heichips25_sap3/_0684_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3072_  (.B1(\heichips25_sap3/_1548_ ),
    .Y(\heichips25_sap3/_0685_ ),
    .A1(\heichips25_sap3/_1464_ ),
    .A2(\heichips25_sap3/_1552_ ));
 sg13g2_nand3_1 \heichips25_sap3/_3073_  (.B(\heichips25_sap3/net245 ),
    .C(\heichips25_sap3/_0685_ ),
    .A(\heichips25_sap3/net266 ),
    .Y(\heichips25_sap3/_0686_ ));
 sg13g2_nor3_1 \heichips25_sap3/_3074_  (.A(\heichips25_sap3/_1486_ ),
    .B(\heichips25_sap3/_1495_ ),
    .C(\heichips25_sap3/_1508_ ),
    .Y(\heichips25_sap3/_0687_ ));
 sg13g2_a21o_1 \heichips25_sap3/_3075_  (.A2(\heichips25_sap3/_1548_ ),
    .A1(\heichips25_sap3/_1497_ ),
    .B1(\heichips25_sap3/_1518_ ),
    .X(\heichips25_sap3/_0688_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3076_  (.A(\heichips25_sap3/_1462_ ),
    .B(\heichips25_sap3/_1508_ ),
    .Y(\heichips25_sap3/_0689_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_3077_  (.Y(\heichips25_sap3/_0690_ ),
    .B(\heichips25_sap3/net249 ),
    .A_N(\heichips25_sap3/_1668_ ));
 sg13g2_nand3_1 \heichips25_sap3/_3078_  (.B(\heichips25_sap3/_0686_ ),
    .C(\heichips25_sap3/_0688_ ),
    .A(\heichips25_sap3/_0684_ ),
    .Y(\heichips25_sap3/_0691_ ));
 sg13g2_or4_1 \heichips25_sap3/_3079_  (.A(\heichips25_sap3/_1697_ ),
    .B(\heichips25_sap3/_0648_ ),
    .C(\heichips25_sap3/_0683_ ),
    .D(\heichips25_sap3/_0687_ ),
    .X(\heichips25_sap3/_0692_ ));
 sg13g2_nor3_1 \heichips25_sap3/_3080_  (.A(\heichips25_sap3/_0682_ ),
    .B(\heichips25_sap3/_0691_ ),
    .C(\heichips25_sap3/_0692_ ),
    .Y(\heichips25_sap3/_0693_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3081_  (.A1(\heichips25_sap3/net220 ),
    .A2(\heichips25_sap3/_0689_ ),
    .Y(\heichips25_sap3/_0694_ ),
    .B1(\heichips25_sap3/net249 ));
 sg13g2_o21ai_1 \heichips25_sap3/_3082_  (.B1(\heichips25_sap3/_0694_ ),
    .Y(\heichips25_sap3/_0695_ ),
    .A1(\heichips25_sap3/net220 ),
    .A2(\heichips25_sap3/_0693_ ));
 sg13g2_and3_1 \heichips25_sap3/_3083_  (.X(\heichips25_sap3/_0696_ ),
    .A(\heichips25_sap3/_1753_ ),
    .B(\heichips25_sap3/_0690_ ),
    .C(\heichips25_sap3/_0695_ ));
 sg13g2_nand3_1 \heichips25_sap3/_3084_  (.B(\heichips25_sap3/_0690_ ),
    .C(\heichips25_sap3/_0695_ ),
    .A(\heichips25_sap3/_1753_ ),
    .Y(\heichips25_sap3/_0697_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3085_  (.B1(\heichips25_sap3/_0297_ ),
    .Y(\heichips25_sap3/_0698_ ),
    .A1(\heichips25_sap3/_1495_ ),
    .A2(\heichips25_sap3/_1625_ ));
 sg13g2_nor4_1 \heichips25_sap3/_3086_  (.A(\heichips25_sap3/_1525_ ),
    .B(\heichips25_sap3/_1535_ ),
    .C(\heichips25_sap3/_0638_ ),
    .D(\heichips25_sap3/_0698_ ),
    .Y(\heichips25_sap3/_0699_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3087_  (.A(\heichips25_sap3/_1468_ ),
    .B(\heichips25_sap3/_1552_ ),
    .Y(\heichips25_sap3/_0700_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3088_  (.B1(\heichips25_sap3/_0700_ ),
    .Y(\heichips25_sap3/_0701_ ),
    .A1(\heichips25_sap3/net243 ),
    .A2(\heichips25_sap3/_0307_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3089_  (.Y(\heichips25_sap3/_0702_ ),
    .A(\heichips25_sap3/_1560_ ),
    .B(\heichips25_sap3/net222 ));
 sg13g2_o21ai_1 \heichips25_sap3/_3090_  (.B1(\heichips25_sap3/_0307_ ),
    .Y(\heichips25_sap3/_0703_ ),
    .A1(\heichips25_sap3/net236 ),
    .A2(\heichips25_sap3/_0702_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3091_  (.B1(\heichips25_sap3/_0702_ ),
    .Y(\heichips25_sap3/_0704_ ),
    .A1(\heichips25_sap3/net243 ),
    .A2(\heichips25_sap3/_1664_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3092_  (.Y(\heichips25_sap3/_0705_ ),
    .A(\heichips25_sap3/net235 ),
    .B(\heichips25_sap3/net222 ));
 sg13g2_nand4_1 \heichips25_sap3/_3093_  (.B(\heichips25_sap3/_1530_ ),
    .C(\heichips25_sap3/_1544_ ),
    .A(\heichips25_sap3/net271 ),
    .Y(\heichips25_sap3/_0706_ ),
    .D(\heichips25_sap3/_0705_ ));
 sg13g2_and4_1 \heichips25_sap3/_3094_  (.A(\heichips25_sap3/_0701_ ),
    .B(\heichips25_sap3/_0703_ ),
    .C(\heichips25_sap3/_0704_ ),
    .D(\heichips25_sap3/_0706_ ),
    .X(\heichips25_sap3/_0707_ ));
 sg13g2_nor3_1 \heichips25_sap3/_3095_  (.A(\heichips25_sap3/_1503_ ),
    .B(\heichips25_sap3/net242 ),
    .C(\heichips25_sap3/_0295_ ),
    .Y(\heichips25_sap3/_0708_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3096_  (.A(\heichips25_sap3/net222 ),
    .B(\heichips25_sap3/_0708_ ),
    .Y(\heichips25_sap3/_0709_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3097_  (.A1(\heichips25_sap3/_1510_ ),
    .A2(\heichips25_sap3/_0708_ ),
    .Y(\heichips25_sap3/_0710_ ),
    .B1(\heichips25_sap3/net222 ));
 sg13g2_o21ai_1 \heichips25_sap3/_3098_  (.B1(\heichips25_sap3/_1871_ ),
    .Y(\heichips25_sap3/_0711_ ),
    .A1(\heichips25_sap3/net256 ),
    .A2(\heichips25_sap3/_1569_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_3099_  (.B2(\heichips25_sap3/_1526_ ),
    .C1(\heichips25_sap3/_0710_ ),
    .B1(\heichips25_sap3/_0711_ ),
    .A1(\heichips25_sap3/_1524_ ),
    .Y(\heichips25_sap3/_0712_ ),
    .A2(\heichips25_sap3/_1534_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3100_  (.A1(\heichips25_sap3/_0707_ ),
    .A2(\heichips25_sap3/_0712_ ),
    .Y(\heichips25_sap3/_0713_ ),
    .B1(\heichips25_sap3/_0699_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3101_  (.B1(\heichips25_sap3/_0314_ ),
    .Y(\heichips25_sap3/_0714_ ),
    .A1(\heichips25_sap3/_1719_ ),
    .A2(\heichips25_sap3/_0713_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3102_  (.A1(\heichips25_sap3/net247 ),
    .A2(\heichips25_sap3/net246 ),
    .Y(\heichips25_sap3/_0715_ ),
    .B1(\heichips25_sap3/_0654_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3103_  (.Y(\heichips25_sap3/_0716_ ),
    .B1(\heichips25_sap3/_0654_ ),
    .B2(\heichips25_sap3/_1441_ ),
    .A2(\heichips25_sap3/_1467_ ),
    .A1(\heichips25_sap3/_1457_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3104_  (.Y(\heichips25_sap3/_0717_ ),
    .A(\heichips25_sap3/_0714_ ),
    .B(\heichips25_sap3/_0716_ ));
 sg13g2_and3_1 \heichips25_sap3/_3105_  (.X(\heichips25_sap3/_0718_ ),
    .A(\heichips25_sap3/_0697_ ),
    .B(\heichips25_sap3/_0714_ ),
    .C(\heichips25_sap3/_0716_ ));
 sg13g2_and2_1 \heichips25_sap3/_3106_  (.A(\heichips25_sap3/_0680_ ),
    .B(\heichips25_sap3/net152 ),
    .X(\heichips25_sap3/_0719_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3107_  (.Y(\heichips25_sap3/_0720_ ),
    .A(\heichips25_sap3/_0680_ ),
    .B(\heichips25_sap3/net152 ));
 sg13g2_nand2_1 \heichips25_sap3/_3108_  (.Y(\heichips25_sap3/_0721_ ),
    .A(\heichips25_sap3/_0307_ ),
    .B(\heichips25_sap3/_0705_ ));
 sg13g2_nor3_1 \heichips25_sap3/_3109_  (.A(\heichips25_sap3/net242 ),
    .B(\heichips25_sap3/_1664_ ),
    .C(\heichips25_sap3/_0295_ ),
    .Y(\heichips25_sap3/_0722_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3110_  (.A1(\heichips25_sap3/_1513_ ),
    .A2(\heichips25_sap3/_0722_ ),
    .Y(\heichips25_sap3/_0723_ ),
    .B1(\heichips25_sap3/net222 ));
 sg13g2_nor2_1 \heichips25_sap3/_3111_  (.A(\heichips25_sap3/_1565_ ),
    .B(\heichips25_sap3/_1635_ ),
    .Y(\heichips25_sap3/_0724_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3112_  (.A1(\heichips25_sap3/_1504_ ),
    .A2(\heichips25_sap3/_1565_ ),
    .Y(\heichips25_sap3/_0725_ ),
    .B1(\heichips25_sap3/_1480_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3113_  (.B1(\heichips25_sap3/_1509_ ),
    .Y(\heichips25_sap3/_0726_ ),
    .A1(\heichips25_sap3/net230 ),
    .A2(\heichips25_sap3/_1607_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3114_  (.B1(\heichips25_sap3/_0726_ ),
    .Y(\heichips25_sap3/_0727_ ),
    .A1(\heichips25_sap3/_1527_ ),
    .A2(\heichips25_sap3/_1871_ ));
 sg13g2_or4_1 \heichips25_sap3/_3115_  (.A(\heichips25_sap3/_1719_ ),
    .B(\heichips25_sap3/_0698_ ),
    .C(\heichips25_sap3/_0725_ ),
    .D(\heichips25_sap3/_0727_ ),
    .X(\heichips25_sap3/_0728_ ));
 sg13g2_nor3_1 \heichips25_sap3/_3116_  (.A(\heichips25_sap3/_0723_ ),
    .B(\heichips25_sap3/_0724_ ),
    .C(\heichips25_sap3/_0728_ ),
    .Y(\heichips25_sap3/_0729_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3117_  (.A1(\heichips25_sap3/_0721_ ),
    .A2(\heichips25_sap3/_0729_ ),
    .Y(\heichips25_sap3/_0730_ ),
    .B1(\heichips25_sap3/_0313_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_3118_  (.B2(\heichips25_sap3/_1363_ ),
    .C1(\heichips25_sap3/_0730_ ),
    .B1(\heichips25_sap3/_0654_ ),
    .A1(\heichips25_sap3/net247 ),
    .Y(\heichips25_sap3/_0731_ ),
    .A2(\heichips25_sap3/net246 ));
 sg13g2_inv_1 \heichips25_sap3/_3119_  (.Y(\heichips25_sap3/_0732_ ),
    .A(\heichips25_sap3/_0731_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3120_  (.B1(\heichips25_sap3/_1581_ ),
    .Y(\heichips25_sap3/_0733_ ),
    .A1(\heichips25_sap3/net243 ),
    .A2(\heichips25_sap3/_0307_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_3121_  (.B2(\heichips25_sap3/net266 ),
    .C1(\heichips25_sap3/_0724_ ),
    .B1(\heichips25_sap3/_0654_ ),
    .A1(\heichips25_sap3/_1513_ ),
    .Y(\heichips25_sap3/_0734_ ),
    .A2(\heichips25_sap3/_0638_ ));
 sg13g2_or2_1 \heichips25_sap3/_3122_  (.X(\heichips25_sap3/_0735_ ),
    .B(\heichips25_sap3/_1635_ ),
    .A(\heichips25_sap3/_1532_ ));
 sg13g2_nand3_1 \heichips25_sap3/_3123_  (.B(\heichips25_sap3/_0734_ ),
    .C(\heichips25_sap3/_0735_ ),
    .A(\heichips25_sap3/_0733_ ),
    .Y(\heichips25_sap3/_0736_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3124_  (.A(\heichips25_sap3/_0732_ ),
    .B(\heichips25_sap3/net166 ),
    .Y(\heichips25_sap3/_0737_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3125_  (.A1(\heichips25_sap3/_1554_ ),
    .A2(\heichips25_sap3/net225 ),
    .Y(\heichips25_sap3/_0738_ ),
    .B1(\heichips25_sap3/_1536_ ));
 sg13g2_nand4_1 \heichips25_sap3/_3126_  (.B(\heichips25_sap3/_1665_ ),
    .C(\heichips25_sap3/_0646_ ),
    .A(\heichips25_sap3/_1621_ ),
    .Y(\heichips25_sap3/_0739_ ),
    .D(\heichips25_sap3/_0688_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3127_  (.B1(\heichips25_sap3/_1485_ ),
    .Y(\heichips25_sap3/_0740_ ),
    .A1(\heichips25_sap3/_1664_ ),
    .A2(\heichips25_sap3/_0669_ ));
 sg13g2_nand3_1 \heichips25_sap3/_3128_  (.B(\heichips25_sap3/_1758_ ),
    .C(\heichips25_sap3/_0740_ ),
    .A(\heichips25_sap3/_1659_ ),
    .Y(\heichips25_sap3/_0741_ ));
 sg13g2_nor3_1 \heichips25_sap3/_3129_  (.A(\heichips25_sap3/_0738_ ),
    .B(\heichips25_sap3/_0739_ ),
    .C(\heichips25_sap3/_0741_ ),
    .Y(\heichips25_sap3/_0742_ ));
 sg13g2_and2_1 \heichips25_sap3/_3130_  (.A(\heichips25_sap3/_0643_ ),
    .B(\heichips25_sap3/_0742_ ),
    .X(\heichips25_sap3/_0743_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3131_  (.B1(\heichips25_sap3/_0656_ ),
    .Y(\heichips25_sap3/_0744_ ),
    .A1(\heichips25_sap3/_0435_ ),
    .A2(\heichips25_sap3/_0743_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3132_  (.A1(\heichips25_sap3/_1454_ ),
    .A2(\heichips25_sap3/_0744_ ),
    .Y(\heichips25_sap3/_0745_ ),
    .B1(\heichips25_sap3/net249 ));
 sg13g2_nand2b_1 \heichips25_sap3/_3133_  (.Y(\heichips25_sap3/_0746_ ),
    .B(\heichips25_sap3/_0662_ ),
    .A_N(\heichips25_sap3/_0745_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3134_  (.A1(\heichips25_sap3/_0737_ ),
    .A2(\heichips25_sap3/_0746_ ),
    .Y(\heichips25_sap3/_0747_ ),
    .B1(\heichips25_sap3/net123 ));
 sg13g2_inv_1 \heichips25_sap3/_3135_  (.Y(\heichips25_sap3/_0748_ ),
    .A(\heichips25_sap3/_0747_ ));
 sg13g2_and2_1 \heichips25_sap3/_3136_  (.A(\heichips25_sap3/_0731_ ),
    .B(\heichips25_sap3/net166 ),
    .X(\heichips25_sap3/_0749_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3137_  (.Y(\heichips25_sap3/_0750_ ),
    .A(\heichips25_sap3/_0731_ ),
    .B(\heichips25_sap3/net166 ));
 sg13g2_nor2_1 \heichips25_sap3/_3138_  (.A(\heichips25_sap3/_0667_ ),
    .B(\heichips25_sap3/_0679_ ),
    .Y(\heichips25_sap3/_0751_ ));
 sg13g2_and2_1 \heichips25_sap3/_3139_  (.A(\heichips25_sap3/_0717_ ),
    .B(\heichips25_sap3/net151 ),
    .X(\heichips25_sap3/_0752_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3140_  (.Y(\heichips25_sap3/_0753_ ),
    .A(\heichips25_sap3/_0717_ ),
    .B(\heichips25_sap3/net150 ));
 sg13g2_a221oi_1 \heichips25_sap3/_3141_  (.B2(\heichips25_sap3/_0716_ ),
    .C1(\heichips25_sap3/_0679_ ),
    .B1(\heichips25_sap3/_0714_ ),
    .A1(\heichips25_sap3/_0660_ ),
    .Y(\heichips25_sap3/_0754_ ),
    .A2(\heichips25_sap3/_0665_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3142_  (.Y(\heichips25_sap3/_0755_ ),
    .A(\heichips25_sap3/_0680_ ),
    .B(\heichips25_sap3/_0717_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_3143_  (.B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][0] ),
    .C1(\heichips25_sap3/net128 ),
    .B1(\heichips25_sap3/net147 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][0] ),
    .Y(\heichips25_sap3/_0756_ ),
    .A2(\heichips25_sap3/net116 ));
 sg13g2_and2_1 \heichips25_sap3/_3144_  (.A(\heichips25_sap3/net152 ),
    .B(\heichips25_sap3/net150 ),
    .X(\heichips25_sap3/_0757_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3145_  (.Y(\heichips25_sap3/_0758_ ),
    .A(\heichips25_sap3/net152 ),
    .B(\heichips25_sap3/net150 ));
 sg13g2_a221oi_1 \heichips25_sap3/_3146_  (.B2(\heichips25_sap3/_0677_ ),
    .C1(\heichips25_sap3/_0664_ ),
    .B1(\heichips25_sap3/_0676_ ),
    .A1(\heichips25_sap3/net241 ),
    .Y(\heichips25_sap3/_0759_ ),
    .A2(\heichips25_sap3/_0659_ ));
 sg13g2_and4_1 \heichips25_sap3/_3147_  (.A(\heichips25_sap3/_0697_ ),
    .B(\heichips25_sap3/_0714_ ),
    .C(\heichips25_sap3/_0716_ ),
    .D(\heichips25_sap3/_0759_ ),
    .X(\heichips25_sap3/_0760_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3148_  (.Y(\heichips25_sap3/_0761_ ),
    .B1(\heichips25_sap3/net145 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][0] ),
    .A2(\heichips25_sap3/net108 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][0] ));
 sg13g2_nor2_1 \heichips25_sap3/_3149_  (.A(\heichips25_sap3/_0666_ ),
    .B(\heichips25_sap3/_0678_ ),
    .Y(\heichips25_sap3/_0762_ ));
 sg13g2_and2_1 \heichips25_sap3/_3150_  (.A(\heichips25_sap3/net152 ),
    .B(\heichips25_sap3/_0762_ ),
    .X(\heichips25_sap3/_0763_ ));
 sg13g2_inv_1 \heichips25_sap3/_3151_  (.Y(\heichips25_sap3/_0764_ ),
    .A(\heichips25_sap3/net104 ));
 sg13g2_nand2_1 \heichips25_sap3/_3152_  (.Y(\heichips25_sap3/_0765_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][0] ),
    .B(\heichips25_sap3/net105 ));
 sg13g2_nor3_1 \heichips25_sap3/_3153_  (.A(\heichips25_sap3/_0667_ ),
    .B(\heichips25_sap3/_0679_ ),
    .C(\heichips25_sap3/_0697_ ),
    .Y(\heichips25_sap3/_0766_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3154_  (.Y(\heichips25_sap3/_0767_ ),
    .A(\heichips25_sap3/_0696_ ),
    .B(\heichips25_sap3/net150 ));
 sg13g2_nor3_1 \heichips25_sap3/_3155_  (.A(\heichips25_sap3/_0666_ ),
    .B(\heichips25_sap3/_0678_ ),
    .C(\heichips25_sap3/_0697_ ),
    .Y(\heichips25_sap3/_0768_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3156_  (.Y(\heichips25_sap3/_0769_ ),
    .B1(\heichips25_sap3/net138 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][0] ),
    .A2(\heichips25_sap3/net140 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][0] ));
 sg13g2_nor3_1 \heichips25_sap3/_3157_  (.A(\heichips25_sap3/_0666_ ),
    .B(\heichips25_sap3/_0679_ ),
    .C(\heichips25_sap3/_0697_ ),
    .Y(\heichips25_sap3/_0770_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3158_  (.Y(\heichips25_sap3/_0771_ ),
    .A(\heichips25_sap3/_0680_ ),
    .B(\heichips25_sap3/_0696_ ));
 sg13g2_and2_1 \heichips25_sap3/_3159_  (.A(\heichips25_sap3/_0696_ ),
    .B(\heichips25_sap3/_0759_ ),
    .X(\heichips25_sap3/_0772_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3160_  (.Y(\heichips25_sap3/_0773_ ),
    .B1(\heichips25_sap3/net133 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][0] ),
    .A2(\heichips25_sap3/net134 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][0] ));
 sg13g2_and2_1 \heichips25_sap3/_3161_  (.A(\heichips25_sap3/_0769_ ),
    .B(\heichips25_sap3/_0773_ ),
    .X(\heichips25_sap3/_0774_ ));
 sg13g2_nand4_1 \heichips25_sap3/_3162_  (.B(\heichips25_sap3/_0761_ ),
    .C(\heichips25_sap3/_0765_ ),
    .A(\heichips25_sap3/_0756_ ),
    .Y(\heichips25_sap3/_0775_ ),
    .D(\heichips25_sap3/_0774_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3163_  (.Y(\heichips25_sap3/_0776_ ),
    .A(\heichips25_sap3/_1392_ ),
    .B(\heichips25_sap3/net127 ));
 sg13g2_and2_1 \heichips25_sap3/_3164_  (.A(\heichips25_sap3/_0775_ ),
    .B(\heichips25_sap3/_0776_ ),
    .X(\heichips25_sap3/_0777_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3165_  (.Y(\heichips25_sap3/_0778_ ),
    .A(\heichips25_sap3/_0775_ ),
    .B(\heichips25_sap3/_0776_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3166_  (.Y(\heichips25_sap3/_0779_ ),
    .B1(\heichips25_sap3/net147 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][7] ),
    .A2(\heichips25_sap3/net117 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][7] ));
 sg13g2_a22oi_1 \heichips25_sap3/_3167_  (.Y(\heichips25_sap3/_0780_ ),
    .B1(\heichips25_sap3/net135 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][7] ),
    .A2(\heichips25_sap3/net139 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][7] ));
 sg13g2_a22oi_1 \heichips25_sap3/_3168_  (.Y(\heichips25_sap3/_0781_ ),
    .B1(\heichips25_sap3/net132 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][7] ),
    .A2(\heichips25_sap3/net142 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][7] ));
 sg13g2_nand3_1 \heichips25_sap3/_3169_  (.B(\heichips25_sap3/_0780_ ),
    .C(\heichips25_sap3/_0781_ ),
    .A(\heichips25_sap3/_0779_ ),
    .Y(\heichips25_sap3/_0782_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3170_  (.Y(\heichips25_sap3/_0783_ ),
    .B1(\heichips25_sap3/net104 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][7] ),
    .A2(\heichips25_sap3/net109 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][7] ));
 sg13g2_a22oi_1 \heichips25_sap3/_3171_  (.Y(\heichips25_sap3/_0784_ ),
    .B1(\heichips25_sap3/net144 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][7] ),
    .A2(\heichips25_sap3/net128 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][7] ));
 sg13g2_nand2_1 \heichips25_sap3/_3172_  (.Y(\heichips25_sap3/_0785_ ),
    .A(\heichips25_sap3/_0783_ ),
    .B(\heichips25_sap3/_0784_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3173_  (.A(\heichips25_sap3/_0782_ ),
    .B(\heichips25_sap3/_0785_ ),
    .Y(\heichips25_sap3/_0786_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3174_  (.Y(\heichips25_sap3/_0787_ ),
    .B1(\heichips25_sap3/net132 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][6] ),
    .A2(\heichips25_sap3/net139 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][6] ));
 sg13g2_a22oi_1 \heichips25_sap3/_3175_  (.Y(\heichips25_sap3/_0788_ ),
    .B1(\heichips25_sap3/net135 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][6] ),
    .A2(\heichips25_sap3/net142 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][6] ));
 sg13g2_nand2_1 \heichips25_sap3/_3176_  (.Y(\heichips25_sap3/_0789_ ),
    .A(\heichips25_sap3/_0787_ ),
    .B(\heichips25_sap3/_0788_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_3177_  (.B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][6] ),
    .C1(\heichips25_sap3/_0789_ ),
    .B1(\heichips25_sap3/net148 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][6] ),
    .Y(\heichips25_sap3/_0790_ ),
    .A2(\heichips25_sap3/net117 ));
 sg13g2_nand2_1 \heichips25_sap3/_3178_  (.Y(\heichips25_sap3/_0791_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][6] ),
    .B(\heichips25_sap3/net104 ));
 sg13g2_nand2_1 \heichips25_sap3/_3179_  (.Y(\heichips25_sap3/_0792_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][6] ),
    .B(\heichips25_sap3/net144 ));
 sg13g2_a22oi_1 \heichips25_sap3/_3180_  (.Y(\heichips25_sap3/_0793_ ),
    .B1(\heichips25_sap3/net109 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][6] ),
    .A2(\heichips25_sap3/net129 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][6] ));
 sg13g2_and4_1 \heichips25_sap3/_3181_  (.A(\heichips25_sap3/_0790_ ),
    .B(\heichips25_sap3/_0791_ ),
    .C(\heichips25_sap3/_0792_ ),
    .D(\heichips25_sap3/_0793_ ),
    .X(\heichips25_sap3/_0794_ ));
 sg13g2_nand4_1 \heichips25_sap3/_3182_  (.B(\heichips25_sap3/_0791_ ),
    .C(\heichips25_sap3/_0792_ ),
    .A(\heichips25_sap3/_0790_ ),
    .Y(\heichips25_sap3/_0795_ ),
    .D(\heichips25_sap3/_0793_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3183_  (.Y(\heichips25_sap3/_0796_ ),
    .B1(\heichips25_sap3/net148 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][5] ),
    .A2(\heichips25_sap3/net116 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][5] ));
 sg13g2_a22oi_1 \heichips25_sap3/_3184_  (.Y(\heichips25_sap3/_0797_ ),
    .B1(\heichips25_sap3/net132 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][5] ),
    .A2(\heichips25_sap3/net139 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][5] ));
 sg13g2_a22oi_1 \heichips25_sap3/_3185_  (.Y(\heichips25_sap3/_0798_ ),
    .B1(\heichips25_sap3/net135 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][5] ),
    .A2(\heichips25_sap3/net142 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][5] ));
 sg13g2_and2_1 \heichips25_sap3/_3186_  (.A(\heichips25_sap3/_0797_ ),
    .B(\heichips25_sap3/_0798_ ),
    .X(\heichips25_sap3/_0799_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3187_  (.Y(\heichips25_sap3/_0800_ ),
    .B1(\heichips25_sap3/net104 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][5] ),
    .A2(\heichips25_sap3/net109 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][5] ));
 sg13g2_a22oi_1 \heichips25_sap3/_3188_  (.Y(\heichips25_sap3/_0801_ ),
    .B1(\heichips25_sap3/net144 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][5] ),
    .A2(\heichips25_sap3/net129 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][5] ));
 sg13g2_nand4_1 \heichips25_sap3/_3189_  (.B(\heichips25_sap3/_0799_ ),
    .C(\heichips25_sap3/_0800_ ),
    .A(\heichips25_sap3/_0796_ ),
    .Y(\heichips25_sap3/_0802_ ),
    .D(\heichips25_sap3/_0801_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3190_  (.Y(\heichips25_sap3/_0803_ ),
    .B1(\heichips25_sap3/net139 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][4] ),
    .A2(\heichips25_sap3/net142 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][4] ));
 sg13g2_a22oi_1 \heichips25_sap3/_3191_  (.Y(\heichips25_sap3/_0804_ ),
    .B1(\heichips25_sap3/net132 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][4] ),
    .A2(\heichips25_sap3/net135 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][4] ));
 sg13g2_nand2_1 \heichips25_sap3/_3192_  (.Y(\heichips25_sap3/_0805_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][4] ),
    .B(\heichips25_sap3/net148 ));
 sg13g2_nand3_1 \heichips25_sap3/_3193_  (.B(\heichips25_sap3/_0717_ ),
    .C(\heichips25_sap3/net151 ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][4] ),
    .Y(\heichips25_sap3/_0806_ ));
 sg13g2_and4_1 \heichips25_sap3/_3194_  (.A(\heichips25_sap3/_0803_ ),
    .B(\heichips25_sap3/_0804_ ),
    .C(\heichips25_sap3/_0805_ ),
    .D(\heichips25_sap3/_0806_ ),
    .X(\heichips25_sap3/_0807_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3195_  (.Y(\heichips25_sap3/_0808_ ),
    .B1(\heichips25_sap3/net109 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][4] ),
    .A2(\heichips25_sap3/net129 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][4] ));
 sg13g2_a22oi_1 \heichips25_sap3/_3196_  (.Y(\heichips25_sap3/_0809_ ),
    .B1(\heichips25_sap3/net104 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][4] ),
    .A2(\heichips25_sap3/net144 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][4] ));
 sg13g2_nand3_1 \heichips25_sap3/_3197_  (.B(\heichips25_sap3/_0808_ ),
    .C(\heichips25_sap3/_0809_ ),
    .A(\heichips25_sap3/_0807_ ),
    .Y(\heichips25_sap3/_0810_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3198_  (.Y(\heichips25_sap3/_0811_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][3] ),
    .B(\heichips25_sap3/net148 ));
 sg13g2_nand3_1 \heichips25_sap3/_3199_  (.B(\heichips25_sap3/_0717_ ),
    .C(\heichips25_sap3/net151 ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][3] ),
    .Y(\heichips25_sap3/_0812_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3200_  (.Y(\heichips25_sap3/_0813_ ),
    .B1(\heichips25_sap3/net138 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][3] ),
    .A2(\heichips25_sap3/net140 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][3] ));
 sg13g2_a22oi_1 \heichips25_sap3/_3201_  (.Y(\heichips25_sap3/_0814_ ),
    .B1(\heichips25_sap3/net133 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][3] ),
    .A2(\heichips25_sap3/net135 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][3] ));
 sg13g2_and4_1 \heichips25_sap3/_3202_  (.A(\heichips25_sap3/_0811_ ),
    .B(\heichips25_sap3/_0812_ ),
    .C(\heichips25_sap3/_0813_ ),
    .D(\heichips25_sap3/_0814_ ),
    .X(\heichips25_sap3/_0815_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3203_  (.Y(\heichips25_sap3/_0816_ ),
    .B1(\heichips25_sap3/net105 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][3] ),
    .A2(\heichips25_sap3/net108 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][3] ));
 sg13g2_nand2_1 \heichips25_sap3/_3204_  (.Y(\heichips25_sap3/_0817_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][3] ),
    .B(\heichips25_sap3/net144 ));
 sg13g2_nand2_1 \heichips25_sap3/_3205_  (.Y(\heichips25_sap3/_0818_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][3] ),
    .B(\heichips25_sap3/net128 ));
 sg13g2_and4_1 \heichips25_sap3/_3206_  (.A(\heichips25_sap3/_0815_ ),
    .B(\heichips25_sap3/_0816_ ),
    .C(\heichips25_sap3/_0817_ ),
    .D(\heichips25_sap3/_0818_ ),
    .X(\heichips25_sap3/_0819_ ));
 sg13g2_nand4_1 \heichips25_sap3/_3207_  (.B(\heichips25_sap3/_0816_ ),
    .C(\heichips25_sap3/_0817_ ),
    .A(\heichips25_sap3/_0815_ ),
    .Y(\heichips25_sap3/_0820_ ),
    .D(\heichips25_sap3/_0818_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3208_  (.Y(\heichips25_sap3/_0821_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][0] ),
    .B(\heichips25_sap3/net147 ));
 sg13g2_nand3_1 \heichips25_sap3/_3209_  (.B(\heichips25_sap3/_0717_ ),
    .C(\heichips25_sap3/net151 ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][0] ),
    .Y(\heichips25_sap3/_0822_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3210_  (.Y(\heichips25_sap3/_0823_ ),
    .B1(\heichips25_sap3/net138 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][0] ),
    .A2(\heichips25_sap3/net140 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][0] ));
 sg13g2_a22oi_1 \heichips25_sap3/_3211_  (.Y(\heichips25_sap3/_0824_ ),
    .B1(\heichips25_sap3/net133 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][0] ),
    .A2(\heichips25_sap3/net134 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][0] ));
 sg13g2_and4_1 \heichips25_sap3/_3212_  (.A(\heichips25_sap3/_0821_ ),
    .B(\heichips25_sap3/_0822_ ),
    .C(\heichips25_sap3/_0823_ ),
    .D(\heichips25_sap3/_0824_ ),
    .X(\heichips25_sap3/_0825_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3213_  (.Y(\heichips25_sap3/_0826_ ),
    .B1(\heichips25_sap3/net105 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][0] ),
    .A2(\heichips25_sap3/net128 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][0] ));
 sg13g2_nand2_1 \heichips25_sap3/_3214_  (.Y(\heichips25_sap3/_0827_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][0] ),
    .B(\heichips25_sap3/net108 ));
 sg13g2_nand2_1 \heichips25_sap3/_3215_  (.Y(\heichips25_sap3/_0828_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][0] ),
    .B(\heichips25_sap3/net145 ));
 sg13g2_and4_1 \heichips25_sap3/_3216_  (.A(\heichips25_sap3/_0825_ ),
    .B(\heichips25_sap3/_0826_ ),
    .C(\heichips25_sap3/_0827_ ),
    .D(\heichips25_sap3/_0828_ ),
    .X(\heichips25_sap3/_0829_ ));
 sg13g2_nand4_1 \heichips25_sap3/_3217_  (.B(\heichips25_sap3/_0826_ ),
    .C(\heichips25_sap3/_0827_ ),
    .A(\heichips25_sap3/_0825_ ),
    .Y(\heichips25_sap3/_0830_ ),
    .D(\heichips25_sap3/_0828_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3218_  (.Y(\heichips25_sap3/_0831_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][2] ),
    .B(\heichips25_sap3/net147 ));
 sg13g2_nand3_1 \heichips25_sap3/_3219_  (.B(\heichips25_sap3/_0717_ ),
    .C(\heichips25_sap3/net150 ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][2] ),
    .Y(\heichips25_sap3/_0832_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3220_  (.Y(\heichips25_sap3/_0833_ ),
    .B1(\heichips25_sap3/net138 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][2] ),
    .A2(\heichips25_sap3/net140 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][2] ));
 sg13g2_a22oi_1 \heichips25_sap3/_3221_  (.Y(\heichips25_sap3/_0834_ ),
    .B1(\heichips25_sap3/net133 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][2] ),
    .A2(\heichips25_sap3/net134 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][2] ));
 sg13g2_and4_1 \heichips25_sap3/_3222_  (.A(\heichips25_sap3/_0831_ ),
    .B(\heichips25_sap3/_0832_ ),
    .C(\heichips25_sap3/_0833_ ),
    .D(\heichips25_sap3/_0834_ ),
    .X(\heichips25_sap3/_0835_ ));
 sg13g2_nand3_1 \heichips25_sap3/_3223_  (.B(\heichips25_sap3/net152 ),
    .C(\heichips25_sap3/net150 ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][2] ),
    .Y(\heichips25_sap3/_0836_ ));
 sg13g2_nand3_1 \heichips25_sap3/_3224_  (.B(\heichips25_sap3/net152 ),
    .C(\heichips25_sap3/_0762_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][2] ),
    .Y(\heichips25_sap3/_0837_ ));
 sg13g2_nand3_1 \heichips25_sap3/_3225_  (.B(\heichips25_sap3/_0680_ ),
    .C(\heichips25_sap3/net152 ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][2] ),
    .Y(\heichips25_sap3/_0838_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3226_  (.Y(\heichips25_sap3/_0839_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][2] ),
    .B(\heichips25_sap3/net145 ));
 sg13g2_and4_1 \heichips25_sap3/_3227_  (.A(\heichips25_sap3/_0836_ ),
    .B(\heichips25_sap3/_0837_ ),
    .C(\heichips25_sap3/_0838_ ),
    .D(\heichips25_sap3/_0839_ ),
    .X(\heichips25_sap3/_0840_ ));
 sg13g2_and2_1 \heichips25_sap3/_3228_  (.A(\heichips25_sap3/_0835_ ),
    .B(\heichips25_sap3/_0840_ ),
    .X(\heichips25_sap3/_0841_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3229_  (.Y(\heichips25_sap3/_0842_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][1] ),
    .B(\heichips25_sap3/net147 ));
 sg13g2_nand3_1 \heichips25_sap3/_3230_  (.B(\heichips25_sap3/_0717_ ),
    .C(\heichips25_sap3/net150 ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][1] ),
    .Y(\heichips25_sap3/_0843_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3231_  (.Y(\heichips25_sap3/_0844_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][1] ),
    .B(\heichips25_sap3/net134 ));
 sg13g2_nand3_1 \heichips25_sap3/_3232_  (.B(\heichips25_sap3/_0718_ ),
    .C(\heichips25_sap3/net150 ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][1] ),
    .Y(\heichips25_sap3/_0845_ ));
 sg13g2_nand3_1 \heichips25_sap3/_3233_  (.B(\heichips25_sap3/_0680_ ),
    .C(\heichips25_sap3/_0718_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][1] ),
    .Y(\heichips25_sap3/_0846_ ));
 sg13g2_nand3_1 \heichips25_sap3/_3234_  (.B(\heichips25_sap3/_0718_ ),
    .C(\heichips25_sap3/_0762_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][1] ),
    .Y(\heichips25_sap3/_0847_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3235_  (.Y(\heichips25_sap3/_0848_ ),
    .B1(\heichips25_sap3/net138 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][1] ),
    .A2(\heichips25_sap3/net145 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][1] ));
 sg13g2_a22oi_1 \heichips25_sap3/_3236_  (.Y(\heichips25_sap3/_0849_ ),
    .B1(\heichips25_sap3/net133 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][1] ),
    .A2(\heichips25_sap3/net140 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][1] ));
 sg13g2_and4_1 \heichips25_sap3/_3237_  (.A(\heichips25_sap3/_0844_ ),
    .B(\heichips25_sap3/_0846_ ),
    .C(\heichips25_sap3/_0848_ ),
    .D(\heichips25_sap3/_0849_ ),
    .X(\heichips25_sap3/_0850_ ));
 sg13g2_and4_1 \heichips25_sap3/_3238_  (.A(\heichips25_sap3/_0842_ ),
    .B(\heichips25_sap3/_0843_ ),
    .C(\heichips25_sap3/_0845_ ),
    .D(\heichips25_sap3/_0847_ ),
    .X(\heichips25_sap3/_0851_ ));
 sg13g2_and2_1 \heichips25_sap3/_3239_  (.A(\heichips25_sap3/_0850_ ),
    .B(\heichips25_sap3/_0851_ ),
    .X(\heichips25_sap3/_0852_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3240_  (.Y(\heichips25_sap3/_0853_ ),
    .A(\heichips25_sap3/_0841_ ),
    .B(\heichips25_sap3/_0852_ ));
 sg13g2_nand3_1 \heichips25_sap3/_3241_  (.B(\heichips25_sap3/_0841_ ),
    .C(\heichips25_sap3/_0852_ ),
    .A(\heichips25_sap3/net61 ),
    .Y(\heichips25_sap3/_0854_ ));
 sg13g2_nand4_1 \heichips25_sap3/_3242_  (.B(\heichips25_sap3/net61 ),
    .C(\heichips25_sap3/_0841_ ),
    .A(\heichips25_sap3/_0819_ ),
    .Y(\heichips25_sap3/_0855_ ),
    .D(\heichips25_sap3/_0852_ ));
 sg13g2_nor3_1 \heichips25_sap3/_3243_  (.A(\heichips25_sap3/_0802_ ),
    .B(\heichips25_sap3/net63 ),
    .C(\heichips25_sap3/_0855_ ),
    .Y(\heichips25_sap3/_0856_ ));
 sg13g2_nor4_1 \heichips25_sap3/_3244_  (.A(\heichips25_sap3/_0795_ ),
    .B(\heichips25_sap3/_0802_ ),
    .C(\heichips25_sap3/net63 ),
    .D(\heichips25_sap3/_0855_ ),
    .Y(\heichips25_sap3/_0857_ ));
 sg13g2_and2_1 \heichips25_sap3/_3245_  (.A(\heichips25_sap3/net53 ),
    .B(\heichips25_sap3/_0857_ ),
    .X(\heichips25_sap3/_0858_ ));
 sg13g2_nand3_1 \heichips25_sap3/_3246_  (.B(\heichips25_sap3/net53 ),
    .C(\heichips25_sap3/_0857_ ),
    .A(\heichips25_sap3/_0778_ ),
    .Y(\heichips25_sap3/_0859_ ));
 sg13g2_xnor2_1 \heichips25_sap3/_3247_  (.Y(\heichips25_sap3/_0860_ ),
    .A(\heichips25_sap3/_0777_ ),
    .B(\heichips25_sap3/_0858_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3248_  (.Y(\heichips25_sap3/_0861_ ),
    .A(\heichips25_sap3/net122 ),
    .B(\heichips25_sap3/_0860_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3249_  (.A(\heichips25_sap3/_0731_ ),
    .B(\heichips25_sap3/net166 ),
    .Y(\heichips25_sap3/_0862_ ));
 sg13g2_or2_1 \heichips25_sap3/_3250_  (.X(\heichips25_sap3/_0863_ ),
    .B(\heichips25_sap3/net166 ),
    .A(\heichips25_sap3/_0731_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3251_  (.Y(\heichips25_sap3/_0864_ ),
    .B1(\heichips25_sap3/_0850_ ),
    .B2(\heichips25_sap3/_0851_ ),
    .A2(\heichips25_sap3/_0840_ ),
    .A1(\heichips25_sap3/_0835_ ));
 sg13g2_or2_1 \heichips25_sap3/_3252_  (.X(\heichips25_sap3/_0865_ ),
    .B(\heichips25_sap3/_0852_ ),
    .A(\heichips25_sap3/_0841_ ));
 sg13g2_and3_1 \heichips25_sap3/_3253_  (.X(\heichips25_sap3/_0866_ ),
    .A(\heichips25_sap3/net63 ),
    .B(\heichips25_sap3/_0820_ ),
    .C(\heichips25_sap3/_0864_ ));
 sg13g2_nand3_1 \heichips25_sap3/_3254_  (.B(\heichips25_sap3/_0820_ ),
    .C(\heichips25_sap3/_0864_ ),
    .A(\heichips25_sap3/net63 ),
    .Y(\heichips25_sap3/_0867_ ));
 sg13g2_nand4_1 \heichips25_sap3/_3255_  (.B(\heichips25_sap3/net63 ),
    .C(\heichips25_sap3/_0820_ ),
    .A(\heichips25_sap3/_0802_ ),
    .Y(\heichips25_sap3/_0868_ ),
    .D(\heichips25_sap3/_0864_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_3256_  (.Y(\heichips25_sap3/_0869_ ),
    .B(\heichips25_sap3/_0795_ ),
    .A_N(\heichips25_sap3/_0868_ ));
 sg13g2_nor3_1 \heichips25_sap3/_3257_  (.A(\heichips25_sap3/net53 ),
    .B(\heichips25_sap3/_0794_ ),
    .C(\heichips25_sap3/_0868_ ),
    .Y(\heichips25_sap3/_0870_ ));
 sg13g2_nor4_1 \heichips25_sap3/_3258_  (.A(\heichips25_sap3/_0778_ ),
    .B(\heichips25_sap3/net53 ),
    .C(\heichips25_sap3/_0794_ ),
    .D(\heichips25_sap3/_0868_ ),
    .Y(\heichips25_sap3/_0871_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3259_  (.A(\heichips25_sap3/net61 ),
    .B(\heichips25_sap3/_0867_ ),
    .Y(\heichips25_sap3/_0872_ ));
 sg13g2_nor3_1 \heichips25_sap3/_3260_  (.A(\heichips25_sap3/_0794_ ),
    .B(\heichips25_sap3/net61 ),
    .C(\heichips25_sap3/_0868_ ),
    .Y(\heichips25_sap3/_0873_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3261_  (.A1(\heichips25_sap3/net59 ),
    .A2(\heichips25_sap3/_0870_ ),
    .Y(\heichips25_sap3/_0874_ ),
    .B1(\heichips25_sap3/_0777_ ));
 sg13g2_a21o_1 \heichips25_sap3/_3262_  (.A2(\heichips25_sap3/net49 ),
    .A1(\heichips25_sap3/net59 ),
    .B1(\heichips25_sap3/_0874_ ),
    .X(\heichips25_sap3/_0875_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3263_  (.Y(\heichips25_sap3/_0876_ ),
    .A(\heichips25_sap3/net98 ),
    .B(\heichips25_sap3/_0875_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3264_  (.B1(\heichips25_sap3/_1573_ ),
    .Y(\heichips25_sap3/_0877_ ),
    .A1(\heichips25_sap3/_1527_ ),
    .A2(\heichips25_sap3/_1569_ ));
 sg13g2_nor4_1 \heichips25_sap3/_3265_  (.A(\heichips25_sap3/_1538_ ),
    .B(\heichips25_sap3/_0709_ ),
    .C(\heichips25_sap3/_0727_ ),
    .D(\heichips25_sap3/_0877_ ),
    .Y(\heichips25_sap3/_0878_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3266_  (.A1(\heichips25_sap3/_0707_ ),
    .A2(\heichips25_sap3/_0878_ ),
    .Y(\heichips25_sap3/_0879_ ),
    .B1(\heichips25_sap3/_0699_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3267_  (.B1(\heichips25_sap3/_0314_ ),
    .Y(\heichips25_sap3/_0880_ ),
    .A1(\heichips25_sap3/_1719_ ),
    .A2(\heichips25_sap3/_0879_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3268_  (.Y(\heichips25_sap3/_0881_ ),
    .A(\heichips25_sap3/_0715_ ),
    .B(\heichips25_sap3/_0880_ ));
 sg13g2_inv_1 \heichips25_sap3/_3269_  (.Y(\heichips25_sap3/_0882_ ),
    .A(\heichips25_sap3/net131 ));
 sg13g2_nor2_1 \heichips25_sap3/_3270_  (.A(\heichips25_sap3/net123 ),
    .B(\heichips25_sap3/_0882_ ),
    .Y(\heichips25_sap3/_0883_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3271_  (.Y(\heichips25_sap3/_0884_ ),
    .A(\heichips25_sap3/net127 ),
    .B(\heichips25_sap3/net131 ));
 sg13g2_nand2_1 \heichips25_sap3/_3272_  (.Y(\heichips25_sap3/_0885_ ),
    .A(\uio_out_sap3[0] ),
    .B(\heichips25_sap3/_0884_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3273_  (.Y(\heichips25_sap3/_0886_ ),
    .A(\uio_oe_sap3[0] ),
    .B(\heichips25_sap3/net68 ));
 sg13g2_nand3_1 \heichips25_sap3/_3274_  (.B(\heichips25_sap3/_0885_ ),
    .C(\heichips25_sap3/_0886_ ),
    .A(\heichips25_sap3/_0737_ ),
    .Y(\heichips25_sap3/_0887_ ));
 sg13g2_nor2b_1 \heichips25_sap3/_3275_  (.A(\heichips25_sap3/_0731_ ),
    .B_N(\heichips25_sap3/net166 ),
    .Y(\heichips25_sap3/_0888_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3276_  (.Y(\heichips25_sap3/_0889_ ),
    .A(\heichips25_sap3/_0732_ ),
    .B(\heichips25_sap3/net166 ));
 sg13g2_nand4_1 \heichips25_sap3/_3277_  (.B(\heichips25_sap3/_0861_ ),
    .C(\heichips25_sap3/_0876_ ),
    .A(\heichips25_sap3/_0747_ ),
    .Y(\heichips25_sap3/_0890_ ),
    .D(\heichips25_sap3/_0887_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3278_  (.B1(\heichips25_sap3/_0890_ ),
    .Y(\heichips25_sap3/_0072_ ),
    .A1(\heichips25_sap3/_1392_ ),
    .A2(\heichips25_sap3/_0747_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3279_  (.Y(\heichips25_sap3/_0891_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[0][1] ),
    .B(\heichips25_sap3/net55 ));
 sg13g2_a22oi_1 \heichips25_sap3/_3280_  (.Y(\heichips25_sap3/_0892_ ),
    .B1(\heichips25_sap3/net134 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][1] ),
    .A2(\heichips25_sap3/net138 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][1] ));
 sg13g2_a22oi_1 \heichips25_sap3/_3281_  (.Y(\heichips25_sap3/_0893_ ),
    .B1(\heichips25_sap3/net145 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][1] ),
    .A2(\heichips25_sap3/net146 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][1] ));
 sg13g2_nand2_1 \heichips25_sap3/_3282_  (.Y(\heichips25_sap3/_0894_ ),
    .A(\heichips25_sap3/net123 ),
    .B(\heichips25_sap3/_0893_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_3283_  (.B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][1] ),
    .C1(\heichips25_sap3/_0894_ ),
    .B1(\heichips25_sap3/net105 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][1] ),
    .Y(\heichips25_sap3/_0895_ ),
    .A2(\heichips25_sap3/net108 ));
 sg13g2_o21ai_1 \heichips25_sap3/_3284_  (.B1(\heichips25_sap3/_0892_ ),
    .Y(\heichips25_sap3/_0896_ ),
    .A1(\heichips25_sap3/_1386_ ),
    .A2(\heichips25_sap3/net115 ));
 sg13g2_a221oi_1 \heichips25_sap3/_3285_  (.B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][1] ),
    .C1(\heichips25_sap3/_0896_ ),
    .B1(\heichips25_sap3/net133 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][1] ),
    .Y(\heichips25_sap3/_0897_ ),
    .A2(\heichips25_sap3/net141 ));
 sg13g2_a22oi_1 \heichips25_sap3/_3286_  (.Y(\heichips25_sap3/_0898_ ),
    .B1(\heichips25_sap3/_0895_ ),
    .B2(\heichips25_sap3/_0897_ ),
    .A2(\heichips25_sap3/net128 ),
    .A1(\heichips25_sap3/_1385_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3287_  (.A(\heichips25_sap3/_0777_ ),
    .B(\heichips25_sap3/net51 ),
    .Y(\heichips25_sap3/_0899_ ));
 sg13g2_nand3_1 \heichips25_sap3/_3288_  (.B(\heichips25_sap3/_0857_ ),
    .C(\heichips25_sap3/_0899_ ),
    .A(\heichips25_sap3/net53 ),
    .Y(\heichips25_sap3/_0900_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3289_  (.Y(\heichips25_sap3/_0901_ ),
    .B1(\heichips25_sap3/_0899_ ),
    .B2(\heichips25_sap3/_0858_ ),
    .A2(\heichips25_sap3/net51 ),
    .A1(\heichips25_sap3/_0859_ ));
 sg13g2_and2_1 \heichips25_sap3/_3290_  (.A(\heichips25_sap3/net61 ),
    .B(\heichips25_sap3/_0852_ ),
    .X(\heichips25_sap3/_0902_ ));
 sg13g2_xnor2_1 \heichips25_sap3/_3291_  (.Y(\heichips25_sap3/_0903_ ),
    .A(\heichips25_sap3/net61 ),
    .B(\heichips25_sap3/_0852_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3292_  (.A(\heichips25_sap3/net127 ),
    .B(\heichips25_sap3/_0903_ ),
    .Y(\heichips25_sap3/_0904_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3293_  (.A1(\heichips25_sap3/net127 ),
    .A2(\heichips25_sap3/_0901_ ),
    .Y(\heichips25_sap3/_0905_ ),
    .B1(\heichips25_sap3/_0904_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3294_  (.Y(\heichips25_sap3/_0906_ ),
    .A(\heichips25_sap3/_1922_ ),
    .B(\heichips25_sap3/_0884_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3295_  (.Y(\heichips25_sap3/_0907_ ),
    .A(\heichips25_sap3/_0327_ ),
    .B(\heichips25_sap3/net68 ));
 sg13g2_a221oi_1 \heichips25_sap3/_3296_  (.B2(\heichips25_sap3/_0907_ ),
    .C1(\heichips25_sap3/_0732_ ),
    .B1(\heichips25_sap3/_0906_ ),
    .A1(\heichips25_sap3/net122 ),
    .Y(\heichips25_sap3/_0908_ ),
    .A2(\heichips25_sap3/_0905_ ));
 sg13g2_nand3_1 \heichips25_sap3/_3297_  (.B(\heichips25_sap3/net48 ),
    .C(\heichips25_sap3/net51 ),
    .A(\heichips25_sap3/net59 ),
    .Y(\heichips25_sap3/_0909_ ));
 sg13g2_a21o_1 \heichips25_sap3/_3298_  (.A2(\heichips25_sap3/net48 ),
    .A1(\heichips25_sap3/net59 ),
    .B1(\heichips25_sap3/net51 ),
    .X(\heichips25_sap3/_0910_ ));
 sg13g2_and2_1 \heichips25_sap3/_3299_  (.A(\heichips25_sap3/_0909_ ),
    .B(\heichips25_sap3/_0910_ ),
    .X(\heichips25_sap3/_0911_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3300_  (.A1(\heichips25_sap3/net127 ),
    .A2(\heichips25_sap3/_0911_ ),
    .Y(\heichips25_sap3/_0912_ ),
    .B1(\heichips25_sap3/_0863_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_3301_  (.Y(\heichips25_sap3/_0913_ ),
    .B(\heichips25_sap3/_0747_ ),
    .A_N(\heichips25_sap3/_0912_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3302_  (.B1(\heichips25_sap3/_0891_ ),
    .Y(\heichips25_sap3/_0073_ ),
    .A1(\heichips25_sap3/_0908_ ),
    .A2(\heichips25_sap3/_0913_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3303_  (.B1(\heichips25_sap3/_0854_ ),
    .Y(\heichips25_sap3/_0914_ ),
    .A1(\heichips25_sap3/_0841_ ),
    .A2(\heichips25_sap3/_0902_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_3304_  (.B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][2] ),
    .C1(\heichips25_sap3/net128 ),
    .B1(\heichips25_sap3/net147 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][2] ),
    .Y(\heichips25_sap3/_0915_ ),
    .A2(\heichips25_sap3/net116 ));
 sg13g2_nand2_1 \heichips25_sap3/_3305_  (.Y(\heichips25_sap3/_0916_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][2] ),
    .B(\heichips25_sap3/net145 ));
 sg13g2_a22oi_1 \heichips25_sap3/_3306_  (.Y(\heichips25_sap3/_0917_ ),
    .B1(\heichips25_sap3/net133 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][2] ),
    .A2(\heichips25_sap3/net140 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][2] ));
 sg13g2_a22oi_1 \heichips25_sap3/_3307_  (.Y(\heichips25_sap3/_0918_ ),
    .B1(\heichips25_sap3/net137 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][2] ),
    .A2(\heichips25_sap3/net138 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][2] ));
 sg13g2_and2_1 \heichips25_sap3/_3308_  (.A(\heichips25_sap3/_0917_ ),
    .B(\heichips25_sap3/_0918_ ),
    .X(\heichips25_sap3/_0919_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3309_  (.Y(\heichips25_sap3/_0920_ ),
    .B1(\heichips25_sap3/net105 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][2] ),
    .A2(\heichips25_sap3/net108 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][2] ));
 sg13g2_and4_1 \heichips25_sap3/_3310_  (.A(\heichips25_sap3/_0915_ ),
    .B(\heichips25_sap3/_0916_ ),
    .C(\heichips25_sap3/_0919_ ),
    .D(\heichips25_sap3/_0920_ ),
    .X(\heichips25_sap3/_0921_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3311_  (.A1(\heichips25_sap3/_1375_ ),
    .A2(\heichips25_sap3/net127 ),
    .Y(\heichips25_sap3/_0922_ ),
    .B1(\heichips25_sap3/_0921_ ));
 sg13g2_xor2_1 \heichips25_sap3/_3312_  (.B(\heichips25_sap3/net50 ),
    .A(\heichips25_sap3/_0900_ ),
    .X(\heichips25_sap3/_0923_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3313_  (.A(\heichips25_sap3/net119 ),
    .B(\heichips25_sap3/_0923_ ),
    .Y(\heichips25_sap3/_0924_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3314_  (.B1(\heichips25_sap3/_0924_ ),
    .Y(\heichips25_sap3/_0925_ ),
    .A1(\heichips25_sap3/net127 ),
    .A2(\heichips25_sap3/_0914_ ));
 sg13g2_nand4_1 \heichips25_sap3/_3315_  (.B(\heichips25_sap3/net48 ),
    .C(\heichips25_sap3/net52 ),
    .A(\heichips25_sap3/net59 ),
    .Y(\heichips25_sap3/_0926_ ),
    .D(\heichips25_sap3/net50 ));
 sg13g2_nand3_1 \heichips25_sap3/_3316_  (.B(\heichips25_sap3/net51 ),
    .C(\heichips25_sap3/net50 ),
    .A(\heichips25_sap3/net48 ),
    .Y(\heichips25_sap3/_0927_ ));
 sg13g2_xnor2_1 \heichips25_sap3/_3317_  (.Y(\heichips25_sap3/_0928_ ),
    .A(\heichips25_sap3/_0909_ ),
    .B(\heichips25_sap3/net50 ));
 sg13g2_nand2_1 \heichips25_sap3/_3318_  (.Y(\heichips25_sap3/_0929_ ),
    .A(\heichips25_sap3/net97 ),
    .B(\heichips25_sap3/_0928_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_3319_  (.Y(\heichips25_sap3/_0930_ ),
    .B(\heichips25_sap3/net68 ),
    .A_N(\uio_oe_sap3[2] ));
 sg13g2_o21ai_1 \heichips25_sap3/_3320_  (.B1(\heichips25_sap3/_0930_ ),
    .Y(\heichips25_sap3/_0931_ ),
    .A1(net44),
    .A2(\heichips25_sap3/net68 ));
 sg13g2_and3_1 \heichips25_sap3/_3321_  (.X(\heichips25_sap3/_0932_ ),
    .A(\heichips25_sap3/_0747_ ),
    .B(\heichips25_sap3/_0929_ ),
    .C(\heichips25_sap3/_0931_ ));
 sg13g2_nand3_1 \heichips25_sap3/_3322_  (.B(\heichips25_sap3/_0865_ ),
    .C(\heichips25_sap3/_0888_ ),
    .A(\heichips25_sap3/_0853_ ),
    .Y(\heichips25_sap3/_0933_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3323_  (.A(\heichips25_sap3/net61 ),
    .B(\heichips25_sap3/_0865_ ),
    .Y(\heichips25_sap3/_0934_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3324_  (.B1(\heichips25_sap3/_0841_ ),
    .Y(\heichips25_sap3/_0935_ ),
    .A1(\heichips25_sap3/net61 ),
    .A2(\heichips25_sap3/_0852_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3325_  (.Y(\heichips25_sap3/_0074_ ),
    .B1(\heichips25_sap3/_0925_ ),
    .B2(\heichips25_sap3/_0932_ ),
    .A2(\heichips25_sap3/net55 ),
    .A1(\heichips25_sap3/_1375_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_3326_  (.B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][3] ),
    .C1(\heichips25_sap3/net128 ),
    .B1(\heichips25_sap3/net148 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][3] ),
    .Y(\heichips25_sap3/_0936_ ),
    .A2(\heichips25_sap3/net116 ));
 sg13g2_a22oi_1 \heichips25_sap3/_3327_  (.Y(\heichips25_sap3/_0937_ ),
    .B1(\heichips25_sap3/net144 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][3] ),
    .A2(\heichips25_sap3/net110 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][3] ));
 sg13g2_nand2_1 \heichips25_sap3/_3328_  (.Y(\heichips25_sap3/_0938_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][3] ),
    .B(\heichips25_sap3/net105 ));
 sg13g2_a22oi_1 \heichips25_sap3/_3329_  (.Y(\heichips25_sap3/_0939_ ),
    .B1(\heichips25_sap3/net133 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][3] ),
    .A2(\heichips25_sap3/net137 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][3] ));
 sg13g2_a22oi_1 \heichips25_sap3/_3330_  (.Y(\heichips25_sap3/_0940_ ),
    .B1(\heichips25_sap3/net138 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][3] ),
    .A2(\heichips25_sap3/net140 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][3] ));
 sg13g2_and2_1 \heichips25_sap3/_3331_  (.A(\heichips25_sap3/_0939_ ),
    .B(\heichips25_sap3/_0940_ ),
    .X(\heichips25_sap3/_0941_ ));
 sg13g2_and4_1 \heichips25_sap3/_3332_  (.A(\heichips25_sap3/_0936_ ),
    .B(\heichips25_sap3/_0937_ ),
    .C(\heichips25_sap3/_0938_ ),
    .D(\heichips25_sap3/_0941_ ),
    .X(\heichips25_sap3/_0942_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3333_  (.A1(\heichips25_sap3/_1368_ ),
    .A2(\heichips25_sap3/net127 ),
    .Y(\heichips25_sap3/_0943_ ),
    .B1(\heichips25_sap3/_0942_ ));
 sg13g2_nand4_1 \heichips25_sap3/_3334_  (.B(\heichips25_sap3/net52 ),
    .C(\heichips25_sap3/net50 ),
    .A(\heichips25_sap3/net48 ),
    .Y(\heichips25_sap3/_0944_ ),
    .D(\heichips25_sap3/_0943_ ));
 sg13g2_inv_1 \heichips25_sap3/_3335_  (.Y(\heichips25_sap3/_0945_ ),
    .A(\heichips25_sap3/_0944_ ));
 sg13g2_xnor2_1 \heichips25_sap3/_3336_  (.Y(\heichips25_sap3/_0946_ ),
    .A(\heichips25_sap3/_0926_ ),
    .B(\heichips25_sap3/_0943_ ));
 sg13g2_xnor2_1 \heichips25_sap3/_3337_  (.Y(\heichips25_sap3/_0947_ ),
    .A(\heichips25_sap3/_0819_ ),
    .B(\heichips25_sap3/_0934_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3338_  (.B1(\heichips25_sap3/net98 ),
    .Y(\heichips25_sap3/_0948_ ),
    .A1(\heichips25_sap3/net128 ),
    .A2(\heichips25_sap3/_0947_ ));
 sg13g2_inv_1 \heichips25_sap3/_3339_  (.Y(\heichips25_sap3/_0949_ ),
    .A(\heichips25_sap3/_0948_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3340_  (.B1(\heichips25_sap3/_0949_ ),
    .Y(\heichips25_sap3/_0950_ ),
    .A1(\heichips25_sap3/net123 ),
    .A2(\heichips25_sap3/_0946_ ));
 sg13g2_nor4_1 \heichips25_sap3/_3341_  (.A(\heichips25_sap3/_0777_ ),
    .B(\heichips25_sap3/net52 ),
    .C(\heichips25_sap3/net50 ),
    .D(\heichips25_sap3/_0943_ ),
    .Y(\heichips25_sap3/_0951_ ));
 sg13g2_nand3_1 \heichips25_sap3/_3342_  (.B(\heichips25_sap3/_0857_ ),
    .C(\heichips25_sap3/_0951_ ),
    .A(\heichips25_sap3/net53 ),
    .Y(\heichips25_sap3/_0952_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3343_  (.B1(\heichips25_sap3/_0943_ ),
    .Y(\heichips25_sap3/_0953_ ),
    .A1(\heichips25_sap3/_0900_ ),
    .A2(\heichips25_sap3/net50 ));
 sg13g2_a21oi_1 \heichips25_sap3/_3344_  (.A1(\heichips25_sap3/_0952_ ),
    .A2(\heichips25_sap3/_0953_ ),
    .Y(\heichips25_sap3/_0954_ ),
    .B1(\heichips25_sap3/net120 ));
 sg13g2_nor2_1 \heichips25_sap3/_3345_  (.A(\uio_oe_sap3[3] ),
    .B(\heichips25_sap3/_0884_ ),
    .Y(\heichips25_sap3/_0955_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3346_  (.A1(\heichips25_sap3/net45 ),
    .A2(\heichips25_sap3/_0884_ ),
    .Y(\heichips25_sap3/_0956_ ),
    .B1(\heichips25_sap3/_0955_ ));
 sg13g2_xnor2_1 \heichips25_sap3/_3347_  (.Y(\heichips25_sap3/_0957_ ),
    .A(\heichips25_sap3/_0819_ ),
    .B(\heichips25_sap3/_0854_ ));
 sg13g2_nor3_1 \heichips25_sap3/_3348_  (.A(\heichips25_sap3/net55 ),
    .B(\heichips25_sap3/_0954_ ),
    .C(\heichips25_sap3/_0956_ ),
    .Y(\heichips25_sap3/_0958_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3349_  (.Y(\heichips25_sap3/_0075_ ),
    .B1(\heichips25_sap3/_0950_ ),
    .B2(\heichips25_sap3/_0958_ ),
    .A2(\heichips25_sap3/net55 ),
    .A1(\heichips25_sap3/_1368_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_3350_  (.B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][4] ),
    .C1(\heichips25_sap3/net129 ),
    .B1(\heichips25_sap3/net148 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][4] ),
    .Y(\heichips25_sap3/_0959_ ),
    .A2(\heichips25_sap3/net116 ));
 sg13g2_nand2_1 \heichips25_sap3/_3351_  (.Y(\heichips25_sap3/_0960_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][4] ),
    .B(\heichips25_sap3/net144 ));
 sg13g2_a22oi_1 \heichips25_sap3/_3352_  (.Y(\heichips25_sap3/_0961_ ),
    .B1(\heichips25_sap3/net132 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][4] ),
    .A2(\heichips25_sap3/net142 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][4] ));
 sg13g2_a22oi_1 \heichips25_sap3/_3353_  (.Y(\heichips25_sap3/_0962_ ),
    .B1(\heichips25_sap3/net135 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][4] ),
    .A2(\heichips25_sap3/net139 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][4] ));
 sg13g2_nand3_1 \heichips25_sap3/_3354_  (.B(\heichips25_sap3/_0961_ ),
    .C(\heichips25_sap3/_0962_ ),
    .A(\heichips25_sap3/_0960_ ),
    .Y(\heichips25_sap3/_0963_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_3355_  (.B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][4] ),
    .C1(\heichips25_sap3/_0963_ ),
    .B1(\heichips25_sap3/net104 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][4] ),
    .Y(\heichips25_sap3/_0964_ ),
    .A2(\heichips25_sap3/net109 ));
 sg13g2_a22oi_1 \heichips25_sap3/_3356_  (.Y(\heichips25_sap3/_0965_ ),
    .B1(\heichips25_sap3/_0959_ ),
    .B2(\heichips25_sap3/_0964_ ),
    .A2(\heichips25_sap3/net129 ),
    .A1(\heichips25_sap3/_1400_ ));
 sg13g2_inv_1 \heichips25_sap3/_3357_  (.Y(\heichips25_sap3/_0966_ ),
    .A(\heichips25_sap3/_0965_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3358_  (.B1(\heichips25_sap3/_0966_ ),
    .Y(\heichips25_sap3/_0967_ ),
    .A1(\heichips25_sap3/net62 ),
    .A2(\heichips25_sap3/_0944_ ));
 sg13g2_and2_1 \heichips25_sap3/_3359_  (.A(\heichips25_sap3/_0943_ ),
    .B(\heichips25_sap3/_0965_ ),
    .X(\heichips25_sap3/_0968_ ));
 sg13g2_nand4_1 \heichips25_sap3/_3360_  (.B(\heichips25_sap3/net52 ),
    .C(\heichips25_sap3/_0922_ ),
    .A(\heichips25_sap3/net49 ),
    .Y(\heichips25_sap3/_0969_ ),
    .D(\heichips25_sap3/_0968_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_3361_  (.Y(\heichips25_sap3/_0970_ ),
    .B(\heichips25_sap3/net59 ),
    .A_N(\heichips25_sap3/_0969_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3362_  (.Y(\heichips25_sap3/_0971_ ),
    .A(\heichips25_sap3/_0967_ ),
    .B(\heichips25_sap3/_0970_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3363_  (.A1(\heichips25_sap3/_0820_ ),
    .A2(\heichips25_sap3/_0934_ ),
    .Y(\heichips25_sap3/_0972_ ),
    .B1(\heichips25_sap3/net63 ));
 sg13g2_nor2_1 \heichips25_sap3/_3364_  (.A(\heichips25_sap3/_0872_ ),
    .B(\heichips25_sap3/_0972_ ),
    .Y(\heichips25_sap3/_0973_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3365_  (.B1(\heichips25_sap3/net96 ),
    .Y(\heichips25_sap3/_0974_ ),
    .A1(\heichips25_sap3/net124 ),
    .A2(\heichips25_sap3/_0973_ ));
 sg13g2_a21o_1 \heichips25_sap3/_3366_  (.A2(\heichips25_sap3/_0971_ ),
    .A1(\heichips25_sap3/net124 ),
    .B1(\heichips25_sap3/_0974_ ),
    .X(\heichips25_sap3/_0975_ ));
 sg13g2_nand4_1 \heichips25_sap3/_3367_  (.B(\heichips25_sap3/_0857_ ),
    .C(\heichips25_sap3/_0951_ ),
    .A(\heichips25_sap3/net53 ),
    .Y(\heichips25_sap3/_0976_ ),
    .D(\heichips25_sap3/_0966_ ));
 sg13g2_xnor2_1 \heichips25_sap3/_3368_  (.Y(\heichips25_sap3/_0977_ ),
    .A(\heichips25_sap3/_0952_ ),
    .B(\heichips25_sap3/_0966_ ));
 sg13g2_xnor2_1 \heichips25_sap3/_3369_  (.Y(\heichips25_sap3/_0978_ ),
    .A(\heichips25_sap3/net63 ),
    .B(\heichips25_sap3/_0855_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3370_  (.B1(\heichips25_sap3/net121 ),
    .Y(\heichips25_sap3/_0979_ ),
    .A1(\heichips25_sap3/net124 ),
    .A2(\heichips25_sap3/_0978_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3371_  (.A1(\heichips25_sap3/net124 ),
    .A2(\heichips25_sap3/_0977_ ),
    .Y(\heichips25_sap3/_0980_ ),
    .B1(\heichips25_sap3/_0979_ ));
 sg13g2_mux2_1 \heichips25_sap3/_3372_  (.A0(net46),
    .A1(\uio_oe_sap3[4] ),
    .S(\heichips25_sap3/net68 ),
    .X(\heichips25_sap3/_0981_ ));
 sg13g2_nor3_1 \heichips25_sap3/_3373_  (.A(\heichips25_sap3/net55 ),
    .B(\heichips25_sap3/_0980_ ),
    .C(\heichips25_sap3/_0981_ ),
    .Y(\heichips25_sap3/_0982_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3374_  (.A1(\heichips25_sap3/_0820_ ),
    .A2(\heichips25_sap3/_0864_ ),
    .Y(\heichips25_sap3/_0983_ ),
    .B1(\heichips25_sap3/_0810_ ));
 sg13g2_nor3_1 \heichips25_sap3/_3375_  (.A(\heichips25_sap3/_0866_ ),
    .B(\heichips25_sap3/_0889_ ),
    .C(\heichips25_sap3/_0983_ ),
    .Y(\heichips25_sap3/_0984_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3376_  (.Y(\heichips25_sap3/_0076_ ),
    .B1(\heichips25_sap3/_0975_ ),
    .B2(\heichips25_sap3/_0982_ ),
    .A2(\heichips25_sap3/net55 ),
    .A1(\heichips25_sap3/_1400_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_3377_  (.B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][5] ),
    .C1(\heichips25_sap3/net124 ),
    .B1(\heichips25_sap3/net146 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][5] ),
    .Y(\heichips25_sap3/_0985_ ),
    .A2(\heichips25_sap3/net116 ));
 sg13g2_nand2_1 \heichips25_sap3/_3378_  (.Y(\heichips25_sap3/_0986_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][5] ),
    .B(\heichips25_sap3/net110 ));
 sg13g2_a22oi_1 \heichips25_sap3/_3379_  (.Y(\heichips25_sap3/_0987_ ),
    .B1(\heichips25_sap3/net139 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][5] ),
    .A2(\heichips25_sap3/net143 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][5] ));
 sg13g2_a22oi_1 \heichips25_sap3/_3380_  (.Y(\heichips25_sap3/_0988_ ),
    .B1(\heichips25_sap3/net132 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][5] ),
    .A2(\heichips25_sap3/net135 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][5] ));
 sg13g2_a22oi_1 \heichips25_sap3/_3381_  (.Y(\heichips25_sap3/_0989_ ),
    .B1(\heichips25_sap3/net104 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][5] ),
    .A2(\heichips25_sap3/_0760_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][5] ));
 sg13g2_and4_1 \heichips25_sap3/_3382_  (.A(\heichips25_sap3/_0986_ ),
    .B(\heichips25_sap3/_0987_ ),
    .C(\heichips25_sap3/_0988_ ),
    .D(\heichips25_sap3/_0989_ ),
    .X(\heichips25_sap3/_0990_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3383_  (.Y(\heichips25_sap3/_0991_ ),
    .B1(\heichips25_sap3/_0985_ ),
    .B2(\heichips25_sap3/_0990_ ),
    .A2(\heichips25_sap3/net124 ),
    .A1(\heichips25_sap3/_1404_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_3384_  (.Y(\heichips25_sap3/_0992_ ),
    .B(\heichips25_sap3/_0991_ ),
    .A_N(\heichips25_sap3/_0969_ ));
 sg13g2_nand3b_1 \heichips25_sap3/_3385_  (.B(\heichips25_sap3/_0991_ ),
    .C(\heichips25_sap3/net59 ),
    .Y(\heichips25_sap3/_0993_ ),
    .A_N(\heichips25_sap3/_0969_ ));
 sg13g2_xnor2_1 \heichips25_sap3/_3386_  (.Y(\heichips25_sap3/_0994_ ),
    .A(\heichips25_sap3/_0970_ ),
    .B(\heichips25_sap3/_0991_ ));
 sg13g2_xnor2_1 \heichips25_sap3/_3387_  (.Y(\heichips25_sap3/_0995_ ),
    .A(\heichips25_sap3/_0802_ ),
    .B(\heichips25_sap3/_0872_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3388_  (.A1(\heichips25_sap3/net123 ),
    .A2(\heichips25_sap3/_0995_ ),
    .Y(\heichips25_sap3/_0996_ ),
    .B1(\heichips25_sap3/_0863_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3389_  (.B1(\heichips25_sap3/_0996_ ),
    .Y(\heichips25_sap3/_0997_ ),
    .A1(\heichips25_sap3/net123 ),
    .A2(\heichips25_sap3/_0994_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3390_  (.A(\heichips25_sap3/_0965_ ),
    .B(\heichips25_sap3/_0991_ ),
    .Y(\heichips25_sap3/_0998_ ));
 sg13g2_and4_1 \heichips25_sap3/_3391_  (.A(\heichips25_sap3/net53 ),
    .B(\heichips25_sap3/_0857_ ),
    .C(\heichips25_sap3/_0951_ ),
    .D(\heichips25_sap3/_0998_ ),
    .X(\heichips25_sap3/_0999_ ));
 sg13g2_nand4_1 \heichips25_sap3/_3392_  (.B(\heichips25_sap3/_0857_ ),
    .C(\heichips25_sap3/_0951_ ),
    .A(\heichips25_sap3/net54 ),
    .Y(\heichips25_sap3/_1000_ ),
    .D(\heichips25_sap3/_0998_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3393_  (.A1(\heichips25_sap3/_0976_ ),
    .A2(\heichips25_sap3/_0991_ ),
    .Y(\heichips25_sap3/_1001_ ),
    .B1(\heichips25_sap3/_0999_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3394_  (.B1(\heichips25_sap3/_0802_ ),
    .Y(\heichips25_sap3/_1002_ ),
    .A1(\heichips25_sap3/net63 ),
    .A2(\heichips25_sap3/_0855_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_3395_  (.Y(\heichips25_sap3/_1003_ ),
    .B(\heichips25_sap3/_1002_ ),
    .A_N(\heichips25_sap3/_0856_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3396_  (.B1(\heichips25_sap3/net121 ),
    .Y(\heichips25_sap3/_1004_ ),
    .A1(\heichips25_sap3/net126 ),
    .A2(\heichips25_sap3/_1003_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3397_  (.A1(\heichips25_sap3/net124 ),
    .A2(\heichips25_sap3/_1001_ ),
    .Y(\heichips25_sap3/_1005_ ),
    .B1(\heichips25_sap3/_1004_ ));
 sg13g2_mux2_1 \heichips25_sap3/_3398_  (.A0(\uio_out_sap3[5] ),
    .A1(\heichips25_sap3/net828 ),
    .S(\heichips25_sap3/net68 ),
    .X(\heichips25_sap3/_1006_ ));
 sg13g2_nor3_1 \heichips25_sap3/_3399_  (.A(\heichips25_sap3/net55 ),
    .B(\heichips25_sap3/_1005_ ),
    .C(\heichips25_sap3/_1006_ ),
    .Y(\heichips25_sap3/_1007_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3400_  (.Y(\heichips25_sap3/_0077_ ),
    .B1(\heichips25_sap3/_0997_ ),
    .B2(\heichips25_sap3/_1007_ ),
    .A2(\heichips25_sap3/net55 ),
    .A1(\heichips25_sap3/_1404_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_3401_  (.B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][6] ),
    .C1(\heichips25_sap3/net126 ),
    .B1(\heichips25_sap3/net146 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][6] ),
    .Y(\heichips25_sap3/_1008_ ),
    .A2(\heichips25_sap3/net116 ));
 sg13g2_nand2_1 \heichips25_sap3/_3402_  (.Y(\heichips25_sap3/_1009_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][6] ),
    .B(\heichips25_sap3/_0763_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3403_  (.Y(\heichips25_sap3/_1010_ ),
    .B1(\heichips25_sap3/net132 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][6] ),
    .A2(\heichips25_sap3/net136 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][6] ));
 sg13g2_a22oi_1 \heichips25_sap3/_3404_  (.Y(\heichips25_sap3/_1011_ ),
    .B1(\heichips25_sap3/_0768_ ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][6] ),
    .A2(\heichips25_sap3/net143 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][6] ));
 sg13g2_nand3_1 \heichips25_sap3/_3405_  (.B(\heichips25_sap3/_1010_ ),
    .C(\heichips25_sap3/_1011_ ),
    .A(\heichips25_sap3/_1009_ ),
    .Y(\heichips25_sap3/_1012_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_3406_  (.B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][6] ),
    .C1(\heichips25_sap3/_1012_ ),
    .B1(\heichips25_sap3/_0760_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][6] ),
    .Y(\heichips25_sap3/_1013_ ),
    .A2(\heichips25_sap3/net110 ));
 sg13g2_a22oi_1 \heichips25_sap3/_3407_  (.Y(\heichips25_sap3/_1014_ ),
    .B1(\heichips25_sap3/_1008_ ),
    .B2(\heichips25_sap3/_1013_ ),
    .A2(\heichips25_sap3/net126 ),
    .A1(\heichips25_sap3/_1412_ ));
 sg13g2_inv_1 \heichips25_sap3/_3408_  (.Y(\heichips25_sap3/_1015_ ),
    .A(\heichips25_sap3/_1014_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3409_  (.Y(\heichips25_sap3/_1016_ ),
    .A(\heichips25_sap3/_0991_ ),
    .B(\heichips25_sap3/_1014_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3410_  (.A(\heichips25_sap3/_0969_ ),
    .B(\heichips25_sap3/_1016_ ),
    .Y(\heichips25_sap3/_1017_ ));
 sg13g2_nor3_1 \heichips25_sap3/_3411_  (.A(\heichips25_sap3/net62 ),
    .B(\heichips25_sap3/_0969_ ),
    .C(\heichips25_sap3/_1016_ ),
    .Y(\heichips25_sap3/_1018_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3412_  (.A1(\heichips25_sap3/_0993_ ),
    .A2(\heichips25_sap3/_1015_ ),
    .Y(\heichips25_sap3/_1019_ ),
    .B1(\heichips25_sap3/_1018_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3413_  (.B1(\heichips25_sap3/_0794_ ),
    .Y(\heichips25_sap3/_1020_ ),
    .A1(\heichips25_sap3/net62 ),
    .A2(\heichips25_sap3/_0868_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_3414_  (.Y(\heichips25_sap3/_1021_ ),
    .B(\heichips25_sap3/_1020_ ),
    .A_N(\heichips25_sap3/_0873_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3415_  (.A1(\heichips25_sap3/net123 ),
    .A2(\heichips25_sap3/_1021_ ),
    .Y(\heichips25_sap3/_1022_ ),
    .B1(\heichips25_sap3/_0863_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3416_  (.B1(\heichips25_sap3/_1022_ ),
    .Y(\heichips25_sap3/_1023_ ),
    .A1(\heichips25_sap3/net123 ),
    .A2(\heichips25_sap3/_1019_ ));
 sg13g2_xnor2_1 \heichips25_sap3/_3417_  (.Y(\heichips25_sap3/_1024_ ),
    .A(\heichips25_sap3/_0999_ ),
    .B(\heichips25_sap3/_1014_ ));
 sg13g2_xnor2_1 \heichips25_sap3/_3418_  (.Y(\heichips25_sap3/_1025_ ),
    .A(\heichips25_sap3/_0794_ ),
    .B(\heichips25_sap3/_0856_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3419_  (.B1(\heichips25_sap3/net121 ),
    .Y(\heichips25_sap3/_1026_ ),
    .A1(\heichips25_sap3/net126 ),
    .A2(\heichips25_sap3/_1025_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3420_  (.A1(\heichips25_sap3/net126 ),
    .A2(\heichips25_sap3/_1024_ ),
    .Y(\heichips25_sap3/_1027_ ),
    .B1(\heichips25_sap3/_1026_ ));
 sg13g2_mux2_1 \heichips25_sap3/_3421_  (.A0(net43),
    .A1(\uio_oe_sap3[6] ),
    .S(\heichips25_sap3/net68 ),
    .X(\heichips25_sap3/_1028_ ));
 sg13g2_nor3_1 \heichips25_sap3/_3422_  (.A(\heichips25_sap3/_0748_ ),
    .B(\heichips25_sap3/_1027_ ),
    .C(\heichips25_sap3/_1028_ ),
    .Y(\heichips25_sap3/_1029_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3423_  (.Y(\heichips25_sap3/_0078_ ),
    .B1(\heichips25_sap3/_1023_ ),
    .B2(\heichips25_sap3/_1029_ ),
    .A2(\heichips25_sap3/_0748_ ),
    .A1(\heichips25_sap3/_1412_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_3424_  (.B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][7] ),
    .C1(\heichips25_sap3/net124 ),
    .B1(\heichips25_sap3/net146 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][7] ),
    .Y(\heichips25_sap3/_1030_ ),
    .A2(\heichips25_sap3/net118 ));
 sg13g2_a22oi_1 \heichips25_sap3/_3425_  (.Y(\heichips25_sap3/_1031_ ),
    .B1(\heichips25_sap3/net104 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][7] ),
    .A2(\heichips25_sap3/net110 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][7] ));
 sg13g2_nand2_1 \heichips25_sap3/_3426_  (.Y(\heichips25_sap3/_1032_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][7] ),
    .B(\heichips25_sap3/net145 ));
 sg13g2_a22oi_1 \heichips25_sap3/_3427_  (.Y(\heichips25_sap3/_1033_ ),
    .B1(\heichips25_sap3/_0772_ ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][7] ),
    .A2(\heichips25_sap3/net142 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][7] ));
 sg13g2_a22oi_1 \heichips25_sap3/_3428_  (.Y(\heichips25_sap3/_1034_ ),
    .B1(\heichips25_sap3/net136 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][7] ),
    .A2(\heichips25_sap3/_0768_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][7] ));
 sg13g2_and4_1 \heichips25_sap3/_3429_  (.A(\heichips25_sap3/_1031_ ),
    .B(\heichips25_sap3/_1032_ ),
    .C(\heichips25_sap3/_1033_ ),
    .D(\heichips25_sap3/_1034_ ),
    .X(\heichips25_sap3/_1035_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3430_  (.Y(\heichips25_sap3/_1036_ ),
    .B1(\heichips25_sap3/_1030_ ),
    .B2(\heichips25_sap3/_1035_ ),
    .A2(\heichips25_sap3/net125 ),
    .A1(\heichips25_sap3/_1420_ ));
 sg13g2_xor2_1 \heichips25_sap3/_3431_  (.B(\heichips25_sap3/_1036_ ),
    .A(\heichips25_sap3/_1018_ ),
    .X(\heichips25_sap3/_1037_ ));
 sg13g2_xnor2_1 \heichips25_sap3/_3432_  (.Y(\heichips25_sap3/_1038_ ),
    .A(\heichips25_sap3/net54 ),
    .B(\heichips25_sap3/_0873_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3433_  (.B1(\heichips25_sap3/net96 ),
    .Y(\heichips25_sap3/_1039_ ),
    .A1(\heichips25_sap3/net125 ),
    .A2(\heichips25_sap3/_1038_ ));
 sg13g2_inv_1 \heichips25_sap3/_3434_  (.Y(\heichips25_sap3/_1040_ ),
    .A(\heichips25_sap3/_1039_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3435_  (.B1(\heichips25_sap3/_1040_ ),
    .Y(\heichips25_sap3/_1041_ ),
    .A1(\heichips25_sap3/_0720_ ),
    .A2(\heichips25_sap3/_1037_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3436_  (.B1(\heichips25_sap3/_1036_ ),
    .Y(\heichips25_sap3/_1042_ ),
    .A1(\heichips25_sap3/_1000_ ),
    .A2(\heichips25_sap3/_1014_ ));
 sg13g2_nand3b_1 \heichips25_sap3/_3437_  (.B(\heichips25_sap3/_0999_ ),
    .C(\heichips25_sap3/_1015_ ),
    .Y(\heichips25_sap3/_1043_ ),
    .A_N(\heichips25_sap3/_1036_ ));
 sg13g2_nand3_1 \heichips25_sap3/_3438_  (.B(\heichips25_sap3/_1042_ ),
    .C(\heichips25_sap3/_1043_ ),
    .A(\heichips25_sap3/net125 ),
    .Y(\heichips25_sap3/_1044_ ));
 sg13g2_xnor2_1 \heichips25_sap3/_3439_  (.Y(\heichips25_sap3/_1045_ ),
    .A(\heichips25_sap3/net54 ),
    .B(\heichips25_sap3/_0857_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3440_  (.B1(\heichips25_sap3/net121 ),
    .Y(\heichips25_sap3/_1046_ ),
    .A1(\heichips25_sap3/net125 ),
    .A2(\heichips25_sap3/_1045_ ));
 sg13g2_inv_1 \heichips25_sap3/_3441_  (.Y(\heichips25_sap3/_1047_ ),
    .A(\heichips25_sap3/_1046_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3442_  (.A(net47),
    .B(\heichips25_sap3/net68 ),
    .Y(\heichips25_sap3/_1048_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3443_  (.A(\uio_oe_sap3[7] ),
    .B(\heichips25_sap3/_0884_ ),
    .Y(\heichips25_sap3/_1049_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3444_  (.B1(\heichips25_sap3/_0747_ ),
    .Y(\heichips25_sap3/_1050_ ),
    .A1(\heichips25_sap3/_1048_ ),
    .A2(\heichips25_sap3/_1049_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3445_  (.A1(\heichips25_sap3/_1044_ ),
    .A2(\heichips25_sap3/_1047_ ),
    .Y(\heichips25_sap3/_1051_ ),
    .B1(\heichips25_sap3/_1050_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3446_  (.Y(\heichips25_sap3/_0079_ ),
    .B1(\heichips25_sap3/_1041_ ),
    .B2(\heichips25_sap3/_1051_ ),
    .A2(\heichips25_sap3/_0748_ ),
    .A1(\heichips25_sap3/_1420_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3447_  (.A(\heichips25_sap3/net105 ),
    .B(\heichips25_sap3/_0883_ ),
    .Y(\heichips25_sap3/_1052_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3448_  (.A(\heichips25_sap3/net119 ),
    .B(\heichips25_sap3/net59 ),
    .Y(\heichips25_sap3/_1053_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3449_  (.Y(\heichips25_sap3/_1054_ ),
    .A(\heichips25_sap3/net122 ),
    .B(\heichips25_sap3/net62 ));
 sg13g2_a21oi_1 \heichips25_sap3/_3450_  (.A1(\heichips25_sap3/_0736_ ),
    .A2(\heichips25_sap3/net62 ),
    .Y(\heichips25_sap3/_1055_ ),
    .B1(\heichips25_sap3/_0731_ ));
 sg13g2_or3_1 \heichips25_sap3/_3451_  (.A(\uio_out_sap3[0] ),
    .B(\heichips25_sap3/_1053_ ),
    .C(\heichips25_sap3/_1055_ ),
    .X(\heichips25_sap3/_1056_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3452_  (.Y(\heichips25_sap3/_1057_ ),
    .A(\heichips25_sap3/net60 ),
    .B(\heichips25_sap3/net99 ));
 sg13g2_nor2b_1 \heichips25_sap3/_3453_  (.A(\heichips25_sap3/net58 ),
    .B_N(\heichips25_sap3/_1057_ ),
    .Y(\heichips25_sap3/_1058_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3454_  (.Y(\heichips25_sap3/_1059_ ),
    .B1(\heichips25_sap3/_1056_ ),
    .B2(\heichips25_sap3/_1058_ ),
    .A2(\heichips25_sap3/net58 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][0] ));
 sg13g2_inv_1 \heichips25_sap3/_3455_  (.Y(\heichips25_sap3/_0080_ ),
    .A(\heichips25_sap3/_1059_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3456_  (.Y(\heichips25_sap3/_1060_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][1] ),
    .B(\heichips25_sap3/net57 ));
 sg13g2_a21o_1 \heichips25_sap3/_3457_  (.A2(\heichips25_sap3/_0903_ ),
    .A1(\heichips25_sap3/net122 ),
    .B1(\uio_out_sap3[1] ),
    .X(\heichips25_sap3/_1061_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3458_  (.A(\heichips25_sap3/_0863_ ),
    .B(\heichips25_sap3/_0903_ ),
    .Y(\heichips25_sap3/_1062_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3459_  (.A(\heichips25_sap3/_1061_ ),
    .B(\heichips25_sap3/_1062_ ),
    .Y(\heichips25_sap3/_1063_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3460_  (.B1(\heichips25_sap3/_1060_ ),
    .Y(\heichips25_sap3/_0081_ ),
    .A1(\heichips25_sap3/net57 ),
    .A2(\heichips25_sap3/_1063_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3461_  (.A1(\heichips25_sap3/net122 ),
    .A2(\heichips25_sap3/_0914_ ),
    .Y(\heichips25_sap3/_1064_ ),
    .B1(net44));
 sg13g2_nand3b_1 \heichips25_sap3/_3462_  (.B(\heichips25_sap3/_0935_ ),
    .C(\heichips25_sap3/net98 ),
    .Y(\heichips25_sap3/_1065_ ),
    .A_N(\heichips25_sap3/_0934_ ));
 sg13g2_nand3_1 \heichips25_sap3/_3463_  (.B(\heichips25_sap3/_1064_ ),
    .C(\heichips25_sap3/_1065_ ),
    .A(\heichips25_sap3/_0933_ ),
    .Y(\heichips25_sap3/_1066_ ));
 sg13g2_mux2_1 \heichips25_sap3/_3464_  (.A0(\heichips25_sap3/_1066_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][2] ),
    .S(\heichips25_sap3/net58 ),
    .X(\heichips25_sap3/_0082_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3465_  (.B1(\heichips25_sap3/net45 ),
    .Y(\heichips25_sap3/_1067_ ),
    .A1(\heichips25_sap3/net119 ),
    .A2(\heichips25_sap3/_0957_ ));
 sg13g2_a21o_1 \heichips25_sap3/_3466_  (.A2(\heichips25_sap3/_0947_ ),
    .A1(\heichips25_sap3/net98 ),
    .B1(\heichips25_sap3/_1067_ ),
    .X(\heichips25_sap3/_1068_ ));
 sg13g2_mux2_1 \heichips25_sap3/_3467_  (.A0(\heichips25_sap3/_1068_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][3] ),
    .S(\heichips25_sap3/net58 ),
    .X(\heichips25_sap3/_0083_ ));
 sg13g2_a21o_1 \heichips25_sap3/_3468_  (.A2(\heichips25_sap3/_0978_ ),
    .A1(\heichips25_sap3/net121 ),
    .B1(net46),
    .X(\heichips25_sap3/_1069_ ));
 sg13g2_nor3_1 \heichips25_sap3/_3469_  (.A(\heichips25_sap3/net98 ),
    .B(\heichips25_sap3/_0984_ ),
    .C(\heichips25_sap3/_1069_ ),
    .Y(\heichips25_sap3/_1070_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3470_  (.A1(\heichips25_sap3/_0764_ ),
    .A2(\heichips25_sap3/_0973_ ),
    .Y(\heichips25_sap3/_1071_ ),
    .B1(\heichips25_sap3/_0863_ ));
 sg13g2_nor3_1 \heichips25_sap3/_3471_  (.A(\heichips25_sap3/net57 ),
    .B(\heichips25_sap3/_1070_ ),
    .C(\heichips25_sap3/_1071_ ),
    .Y(\heichips25_sap3/_1072_ ));
 sg13g2_a21o_1 \heichips25_sap3/_3472_  (.A2(\heichips25_sap3/net57 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][4] ),
    .B1(\heichips25_sap3/_1072_ ),
    .X(\heichips25_sap3/_0084_ ));
 sg13g2_a21o_1 \heichips25_sap3/_3473_  (.A2(\heichips25_sap3/_1003_ ),
    .A1(\heichips25_sap3/net121 ),
    .B1(\uio_out_sap3[5] ),
    .X(\heichips25_sap3/_1073_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3474_  (.A(\heichips25_sap3/_0863_ ),
    .B(\heichips25_sap3/_0995_ ),
    .Y(\heichips25_sap3/_1074_ ));
 sg13g2_nor3_1 \heichips25_sap3/_3475_  (.A(\heichips25_sap3/net57 ),
    .B(\heichips25_sap3/_1073_ ),
    .C(\heichips25_sap3/_1074_ ),
    .Y(\heichips25_sap3/_1075_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3476_  (.A1(\heichips25_sap3/_1411_ ),
    .A2(\heichips25_sap3/net57 ),
    .Y(\heichips25_sap3/_0085_ ),
    .B1(\heichips25_sap3/_1075_ ));
 sg13g2_and2_1 \heichips25_sap3/_3477_  (.A(\heichips25_sap3/net121 ),
    .B(\heichips25_sap3/_1025_ ),
    .X(\heichips25_sap3/_1076_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3478_  (.A(net43),
    .B(\heichips25_sap3/_1076_ ),
    .Y(\heichips25_sap3/_1077_ ));
 sg13g2_or2_1 \heichips25_sap3/_3479_  (.X(\heichips25_sap3/_1078_ ),
    .B(\heichips25_sap3/_1076_ ),
    .A(net43));
 sg13g2_nor2_1 \heichips25_sap3/_3480_  (.A(\heichips25_sap3/_0863_ ),
    .B(\heichips25_sap3/_1021_ ),
    .Y(\heichips25_sap3/_1079_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3481_  (.A(\heichips25_sap3/net57 ),
    .B(\heichips25_sap3/_1079_ ),
    .Y(\heichips25_sap3/_1080_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3482_  (.Y(\heichips25_sap3/_0086_ ),
    .B1(\heichips25_sap3/_1077_ ),
    .B2(\heichips25_sap3/_1080_ ),
    .A2(\heichips25_sap3/net57 ),
    .A1(\heichips25_sap3/_1419_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3483_  (.Y(\heichips25_sap3/_1081_ ),
    .A(\heichips25_sap3/net98 ),
    .B(\heichips25_sap3/_1038_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3484_  (.A1(\heichips25_sap3/net121 ),
    .A2(\heichips25_sap3/_1045_ ),
    .Y(\heichips25_sap3/_1082_ ),
    .B1(net47));
 sg13g2_nand2_1 \heichips25_sap3/_3485_  (.Y(\heichips25_sap3/_1083_ ),
    .A(\heichips25_sap3/_1081_ ),
    .B(\heichips25_sap3/_1082_ ));
 sg13g2_mux2_1 \heichips25_sap3/_3486_  (.A0(\heichips25_sap3/_1083_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][7] ),
    .S(\heichips25_sap3/net58 ),
    .X(\heichips25_sap3/_0087_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3487_  (.Y(\heichips25_sap3/_1084_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][0] ),
    .B(\heichips25_sap3/net106 ));
 sg13g2_nand2_1 \heichips25_sap3/_3488_  (.Y(\heichips25_sap3/_1085_ ),
    .A(\heichips25_sap3/net108 ),
    .B(\heichips25_sap3/_0876_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3489_  (.A(\heichips25_sap3/net119 ),
    .B(\heichips25_sap3/_0860_ ),
    .Y(\heichips25_sap3/_1086_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3490_  (.A(\heichips25_sap3/net106 ),
    .B(\heichips25_sap3/_0882_ ),
    .Y(\heichips25_sap3/_1087_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3491_  (.Y(\heichips25_sap3/_1088_ ),
    .A(\heichips25_sap3/net108 ),
    .B(\heichips25_sap3/net131 ));
 sg13g2_nor2_1 \heichips25_sap3/_3492_  (.A(\uio_oe_sap3[0] ),
    .B(\heichips25_sap3/_1088_ ),
    .Y(\heichips25_sap3/_1089_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3493_  (.A1(\heichips25_sap3/_0212_ ),
    .A2(\heichips25_sap3/_1088_ ),
    .Y(\heichips25_sap3/_1090_ ),
    .B1(\heichips25_sap3/_1089_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3494_  (.A(\heichips25_sap3/net108 ),
    .B(\heichips25_sap3/_1054_ ),
    .Y(\heichips25_sap3/_1091_ ));
 sg13g2_nor4_1 \heichips25_sap3/_3495_  (.A(\heichips25_sap3/_1055_ ),
    .B(\heichips25_sap3/_1086_ ),
    .C(\heichips25_sap3/_1090_ ),
    .D(\heichips25_sap3/_1091_ ),
    .Y(\heichips25_sap3/_1092_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3496_  (.B1(\heichips25_sap3/_1084_ ),
    .Y(\heichips25_sap3/_0088_ ),
    .A1(\heichips25_sap3/_1085_ ),
    .A2(\heichips25_sap3/_1092_ ));
 sg13g2_and2_1 \heichips25_sap3/_3497_  (.A(\heichips25_sap3/net97 ),
    .B(\heichips25_sap3/_0911_ ),
    .X(\heichips25_sap3/_1093_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3498_  (.A(\heichips25_sap3/net119 ),
    .B(\heichips25_sap3/_0901_ ),
    .Y(\heichips25_sap3/_1094_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3499_  (.A(\heichips25_sap3/_1093_ ),
    .B(\heichips25_sap3/_1094_ ),
    .Y(\heichips25_sap3/_1095_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3500_  (.Y(\heichips25_sap3/_1096_ ),
    .A(\heichips25_sap3/_0737_ ),
    .B(\heichips25_sap3/_1088_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3501_  (.A(\uio_out_sap3[1] ),
    .B(\heichips25_sap3/net131 ),
    .Y(\heichips25_sap3/_1097_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3502_  (.A1(\heichips25_sap3/_0327_ ),
    .A2(\heichips25_sap3/_1096_ ),
    .Y(\heichips25_sap3/_1098_ ),
    .B1(\heichips25_sap3/_1097_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3503_  (.A(\heichips25_sap3/net106 ),
    .B(\heichips25_sap3/_1098_ ),
    .Y(\heichips25_sap3/_1099_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3504_  (.Y(\heichips25_sap3/_0089_ ),
    .B1(\heichips25_sap3/_1095_ ),
    .B2(\heichips25_sap3/_1099_ ),
    .A2(\heichips25_sap3/net106 ),
    .A1(\heichips25_sap3/_1391_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3505_  (.Y(\heichips25_sap3/_1100_ ),
    .A(\heichips25_sap3/net122 ),
    .B(\heichips25_sap3/_0923_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3506_  (.Y(\heichips25_sap3/_1101_ ),
    .A(net44),
    .B(\heichips25_sap3/_1088_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3507_  (.A1(\uio_oe_sap3[2] ),
    .A2(\heichips25_sap3/_1087_ ),
    .Y(\heichips25_sap3/_1102_ ),
    .B1(\heichips25_sap3/net122 ));
 sg13g2_nand2_1 \heichips25_sap3/_3508_  (.Y(\heichips25_sap3/_1103_ ),
    .A(\heichips25_sap3/_1101_ ),
    .B(\heichips25_sap3/_1102_ ));
 sg13g2_or2_1 \heichips25_sap3/_3509_  (.X(\heichips25_sap3/_1104_ ),
    .B(\heichips25_sap3/_0914_ ),
    .A(\heichips25_sap3/net119 ));
 sg13g2_a221oi_1 \heichips25_sap3/_3510_  (.B2(\heichips25_sap3/_1103_ ),
    .C1(\heichips25_sap3/net106 ),
    .B1(\heichips25_sap3/_1100_ ),
    .A1(\heichips25_sap3/net97 ),
    .Y(\heichips25_sap3/_1105_ ),
    .A2(\heichips25_sap3/_0928_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3511_  (.A1(\heichips25_sap3/_1380_ ),
    .A2(\heichips25_sap3/net106 ),
    .Y(\heichips25_sap3/_0090_ ),
    .B1(\heichips25_sap3/_1105_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3512_  (.Y(\heichips25_sap3/_1106_ ),
    .A(\heichips25_sap3/net97 ),
    .B(\heichips25_sap3/_0946_ ));
 sg13g2_nor2b_1 \heichips25_sap3/_3513_  (.A(\heichips25_sap3/_0954_ ),
    .B_N(\heichips25_sap3/_1106_ ),
    .Y(\heichips25_sap3/_1107_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3514_  (.Y(\heichips25_sap3/_1108_ ),
    .B1(\heichips25_sap3/_1096_ ),
    .B2(\heichips25_sap3/_0328_ ),
    .A2(\heichips25_sap3/_0882_ ),
    .A1(\heichips25_sap3/net45 ));
 sg13g2_nor2_1 \heichips25_sap3/_3515_  (.A(\heichips25_sap3/net106 ),
    .B(\heichips25_sap3/_1108_ ),
    .Y(\heichips25_sap3/_1109_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3516_  (.Y(\heichips25_sap3/_0091_ ),
    .B1(\heichips25_sap3/_1107_ ),
    .B2(\heichips25_sap3/_1109_ ),
    .A2(\heichips25_sap3/net106 ),
    .A1(\heichips25_sap3/_1373_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3517_  (.A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][4] ),
    .B(\heichips25_sap3/net109 ),
    .Y(\heichips25_sap3/_1110_ ));
 sg13g2_nand3_1 \heichips25_sap3/_3518_  (.B(\heichips25_sap3/_0967_ ),
    .C(\heichips25_sap3/_0970_ ),
    .A(\heichips25_sap3/net96 ),
    .Y(\heichips25_sap3/_1111_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_3519_  (.Y(\heichips25_sap3/_1112_ ),
    .B(\heichips25_sap3/_1087_ ),
    .A_N(\uio_oe_sap3[4] ));
 sg13g2_o21ai_1 \heichips25_sap3/_3520_  (.B1(\heichips25_sap3/_1112_ ),
    .Y(\heichips25_sap3/_1113_ ),
    .A1(net46),
    .A2(\heichips25_sap3/_1087_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_3521_  (.Y(\heichips25_sap3/_1114_ ),
    .B(\heichips25_sap3/_0749_ ),
    .A_N(\heichips25_sap3/_0977_ ));
 sg13g2_nand4_1 \heichips25_sap3/_3522_  (.B(\heichips25_sap3/_1111_ ),
    .C(\heichips25_sap3/_1113_ ),
    .A(\heichips25_sap3/net109 ),
    .Y(\heichips25_sap3/_1115_ ),
    .D(\heichips25_sap3/_1114_ ));
 sg13g2_nor2b_1 \heichips25_sap3/_3523_  (.A(\heichips25_sap3/_1110_ ),
    .B_N(\heichips25_sap3/_1115_ ),
    .Y(\heichips25_sap3/_0092_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3524_  (.A(\heichips25_sap3/net120 ),
    .B(\heichips25_sap3/_1001_ ),
    .Y(\heichips25_sap3/_1116_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3525_  (.A(\uio_out_sap3[5] ),
    .B(\heichips25_sap3/net131 ),
    .Y(\heichips25_sap3/_1117_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3526_  (.B1(\heichips25_sap3/net120 ),
    .Y(\heichips25_sap3/_1118_ ),
    .A1(\heichips25_sap3/net828 ),
    .A2(\heichips25_sap3/_1088_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3527_  (.B1(\heichips25_sap3/net109 ),
    .Y(\heichips25_sap3/_1119_ ),
    .A1(\heichips25_sap3/_1117_ ),
    .A2(\heichips25_sap3/_1118_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3528_  (.A(\heichips25_sap3/_1116_ ),
    .B(\heichips25_sap3/_1119_ ),
    .Y(\heichips25_sap3/_1120_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3529_  (.Y(\heichips25_sap3/_1121_ ),
    .A(\heichips25_sap3/net97 ),
    .B(\heichips25_sap3/_0994_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3530_  (.Y(\heichips25_sap3/_0093_ ),
    .B1(\heichips25_sap3/_1120_ ),
    .B2(\heichips25_sap3/_1121_ ),
    .A2(\heichips25_sap3/net107 ),
    .A1(\heichips25_sap3/_1410_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3531_  (.Y(\heichips25_sap3/_1122_ ),
    .A(\heichips25_sap3/net96 ),
    .B(\heichips25_sap3/_1019_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3532_  (.A(\heichips25_sap3/net120 ),
    .B(\heichips25_sap3/_1024_ ),
    .Y(\heichips25_sap3/_1123_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3533_  (.A1(\heichips25_sap3/net96 ),
    .A2(\heichips25_sap3/_1019_ ),
    .Y(\heichips25_sap3/_1124_ ),
    .B1(\heichips25_sap3/_1123_ ));
 sg13g2_mux2_1 \heichips25_sap3/_3534_  (.A0(net43),
    .A1(\uio_oe_sap3[6] ),
    .S(\heichips25_sap3/_1087_ ),
    .X(\heichips25_sap3/_1125_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3535_  (.A(\heichips25_sap3/net107 ),
    .B(\heichips25_sap3/_1125_ ),
    .Y(\heichips25_sap3/_1126_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3536_  (.Y(\heichips25_sap3/_0094_ ),
    .B1(\heichips25_sap3/_1124_ ),
    .B2(\heichips25_sap3/_1126_ ),
    .A2(\heichips25_sap3/net107 ),
    .A1(\heichips25_sap3/_1418_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_3537_  (.Y(\heichips25_sap3/_1127_ ),
    .B(\heichips25_sap3/_0888_ ),
    .A_N(\heichips25_sap3/_0870_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3538_  (.A1(\heichips25_sap3/net54 ),
    .A2(\heichips25_sap3/_0869_ ),
    .Y(\heichips25_sap3/_1128_ ),
    .B1(\heichips25_sap3/_1127_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3539_  (.Y(\heichips25_sap3/_1129_ ),
    .A(\heichips25_sap3/net96 ),
    .B(\heichips25_sap3/_1037_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3540_  (.A1(\heichips25_sap3/net96 ),
    .A2(\heichips25_sap3/_1037_ ),
    .Y(\heichips25_sap3/_1130_ ),
    .B1(\heichips25_sap3/_1128_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3541_  (.A1(\heichips25_sap3/_1042_ ),
    .A2(\heichips25_sap3/_1043_ ),
    .Y(\heichips25_sap3/_1131_ ),
    .B1(\heichips25_sap3/net120 ));
 sg13g2_mux2_1 \heichips25_sap3/_3542_  (.A0(net47),
    .A1(\uio_oe_sap3[7] ),
    .S(\heichips25_sap3/_1087_ ),
    .X(\heichips25_sap3/_1132_ ));
 sg13g2_nor3_1 \heichips25_sap3/_3543_  (.A(\heichips25_sap3/net107 ),
    .B(\heichips25_sap3/_1131_ ),
    .C(\heichips25_sap3/_1132_ ),
    .Y(\heichips25_sap3/_1133_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3544_  (.Y(\heichips25_sap3/_0095_ ),
    .B1(\heichips25_sap3/_1130_ ),
    .B2(\heichips25_sap3/_1133_ ),
    .A2(\heichips25_sap3/net107 ),
    .A1(\heichips25_sap3/_1425_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_3545_  (.Y(\heichips25_sap3/_1134_ ),
    .B(\heichips25_sap3/_1088_ ),
    .A_N(\heichips25_sap3/net144 ));
 sg13g2_nand3_1 \heichips25_sap3/_3546_  (.B(\heichips25_sap3/_1057_ ),
    .C(\heichips25_sap3/net56 ),
    .A(\heichips25_sap3/_1056_ ),
    .Y(\heichips25_sap3/_1135_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3547_  (.B1(\heichips25_sap3/_1135_ ),
    .Y(\heichips25_sap3/_0096_ ),
    .A1(\heichips25_sap3/_1395_ ),
    .A2(\heichips25_sap3/net56 ));
 sg13g2_o21ai_1 \heichips25_sap3/_3548_  (.B1(\heichips25_sap3/net56 ),
    .Y(\heichips25_sap3/_1136_ ),
    .A1(\heichips25_sap3/_1061_ ),
    .A2(\heichips25_sap3/_1062_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3549_  (.B1(\heichips25_sap3/_1136_ ),
    .Y(\heichips25_sap3/_0097_ ),
    .A1(\heichips25_sap3/_1390_ ),
    .A2(\heichips25_sap3/net56 ));
 sg13g2_mux2_1 \heichips25_sap3/_3550_  (.A0(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][2] ),
    .A1(\heichips25_sap3/_1066_ ),
    .S(\heichips25_sap3/net56 ),
    .X(\heichips25_sap3/_0098_ ));
 sg13g2_mux2_1 \heichips25_sap3/_3551_  (.A0(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][3] ),
    .A1(\heichips25_sap3/_1068_ ),
    .S(\heichips25_sap3/_1134_ ),
    .X(\heichips25_sap3/_0099_ ));
 sg13g2_and2_1 \heichips25_sap3/_3552_  (.A(\heichips25_sap3/net99 ),
    .B(\heichips25_sap3/_0973_ ),
    .X(\heichips25_sap3/_1137_ ));
 sg13g2_or2_1 \heichips25_sap3/_3553_  (.X(\heichips25_sap3/_1138_ ),
    .B(\heichips25_sap3/_1137_ ),
    .A(\heichips25_sap3/_1069_ ));
 sg13g2_mux2_1 \heichips25_sap3/_3554_  (.A0(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][4] ),
    .A1(\heichips25_sap3/_1138_ ),
    .S(\heichips25_sap3/_1134_ ),
    .X(\heichips25_sap3/_0100_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3555_  (.A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][5] ),
    .B(\heichips25_sap3/net56 ),
    .Y(\heichips25_sap3/_1139_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3556_  (.A(\heichips25_sap3/_1073_ ),
    .B(\heichips25_sap3/_1074_ ),
    .Y(\heichips25_sap3/_1140_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3557_  (.A1(\heichips25_sap3/net56 ),
    .A2(\heichips25_sap3/_1140_ ),
    .Y(\heichips25_sap3/_0101_ ),
    .B1(\heichips25_sap3/_1139_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_3558_  (.Y(\heichips25_sap3/_1141_ ),
    .B(\heichips25_sap3/_1077_ ),
    .A_N(\heichips25_sap3/_1079_ ));
 sg13g2_mux2_1 \heichips25_sap3/_3559_  (.A0(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][6] ),
    .A1(\heichips25_sap3/_1141_ ),
    .S(\heichips25_sap3/_1134_ ),
    .X(\heichips25_sap3/_0102_ ));
 sg13g2_mux2_1 \heichips25_sap3/_3560_  (.A0(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][7] ),
    .A1(\heichips25_sap3/_1083_ ),
    .S(\heichips25_sap3/net56 ),
    .X(\heichips25_sap3/_0103_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3561_  (.Y(\heichips25_sap3/_1142_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][0] ),
    .B(\heichips25_sap3/net100 ));
 sg13g2_nand2_1 \heichips25_sap3/_3562_  (.Y(\heichips25_sap3/_1143_ ),
    .A(\heichips25_sap3/net134 ),
    .B(\heichips25_sap3/_0876_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3563_  (.Y(\heichips25_sap3/_1144_ ),
    .A(\heichips25_sap3/net134 ),
    .B(\heichips25_sap3/net131 ));
 sg13g2_nor2_1 \heichips25_sap3/_3564_  (.A(\uio_oe_sap3[0] ),
    .B(\heichips25_sap3/net95 ),
    .Y(\heichips25_sap3/_1145_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3565_  (.A1(\heichips25_sap3/_0212_ ),
    .A2(\heichips25_sap3/net95 ),
    .Y(\heichips25_sap3/_1146_ ),
    .B1(\heichips25_sap3/_1145_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3566_  (.A(\heichips25_sap3/net134 ),
    .B(\heichips25_sap3/_1054_ ),
    .Y(\heichips25_sap3/_1147_ ));
 sg13g2_nor4_1 \heichips25_sap3/_3567_  (.A(\heichips25_sap3/_1055_ ),
    .B(\heichips25_sap3/_1086_ ),
    .C(\heichips25_sap3/_1146_ ),
    .D(\heichips25_sap3/_1147_ ),
    .Y(\heichips25_sap3/_1148_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3568_  (.B1(\heichips25_sap3/_1142_ ),
    .Y(\heichips25_sap3/_0104_ ),
    .A1(\heichips25_sap3/_1143_ ),
    .A2(\heichips25_sap3/_1148_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3569_  (.B1(\heichips25_sap3/net119 ),
    .Y(\heichips25_sap3/_1149_ ),
    .A1(\uio_oe_sap3[1] ),
    .A2(\heichips25_sap3/net95 ));
 sg13g2_nor2_1 \heichips25_sap3/_3570_  (.A(\heichips25_sap3/_1097_ ),
    .B(\heichips25_sap3/_1149_ ),
    .Y(\heichips25_sap3/_1150_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3571_  (.A(\heichips25_sap3/net100 ),
    .B(\heichips25_sap3/_1150_ ),
    .Y(\heichips25_sap3/_1151_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3572_  (.Y(\heichips25_sap3/_0105_ ),
    .B1(\heichips25_sap3/_1095_ ),
    .B2(\heichips25_sap3/_1151_ ),
    .A2(\heichips25_sap3/net100 ),
    .A1(\heichips25_sap3/_1389_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3573_  (.A(net44),
    .B(\heichips25_sap3/net131 ),
    .Y(\heichips25_sap3/_1152_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3574_  (.A(\uio_oe_sap3[2] ),
    .B(\heichips25_sap3/net95 ),
    .Y(\heichips25_sap3/_1153_ ));
 sg13g2_nor3_1 \heichips25_sap3/_3575_  (.A(\heichips25_sap3/net166 ),
    .B(\heichips25_sap3/_1152_ ),
    .C(\heichips25_sap3/_1153_ ),
    .Y(\heichips25_sap3/_1154_ ));
 sg13g2_nor3_1 \heichips25_sap3/_3576_  (.A(\heichips25_sap3/net100 ),
    .B(\heichips25_sap3/_0924_ ),
    .C(\heichips25_sap3/_1154_ ),
    .Y(\heichips25_sap3/_1155_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3577_  (.Y(\heichips25_sap3/_0106_ ),
    .B1(\heichips25_sap3/_0929_ ),
    .B2(\heichips25_sap3/_1155_ ),
    .A2(\heichips25_sap3/net100 ),
    .A1(\heichips25_sap3/_1379_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3578_  (.A(\uio_oe_sap3[3] ),
    .B(\heichips25_sap3/net95 ),
    .Y(\heichips25_sap3/_1156_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3579_  (.A1(\heichips25_sap3/net45 ),
    .A2(\heichips25_sap3/net95 ),
    .Y(\heichips25_sap3/_1157_ ),
    .B1(\heichips25_sap3/_1156_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3580_  (.A(\heichips25_sap3/net100 ),
    .B(\heichips25_sap3/_1157_ ),
    .Y(\heichips25_sap3/_1158_ ));
 sg13g2_xnor2_1 \heichips25_sap3/_3581_  (.Y(\heichips25_sap3/_1159_ ),
    .A(\heichips25_sap3/_0819_ ),
    .B(\heichips25_sap3/_0864_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3582_  (.Y(\heichips25_sap3/_0107_ ),
    .B1(\heichips25_sap3/_1107_ ),
    .B2(\heichips25_sap3/_1158_ ),
    .A2(\heichips25_sap3/net100 ),
    .A1(\heichips25_sap3/_1372_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3583_  (.A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][4] ),
    .B(\heichips25_sap3/net135 ),
    .Y(\heichips25_sap3/_1160_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_3584_  (.Y(\heichips25_sap3/_1161_ ),
    .B(\heichips25_sap3/net95 ),
    .A_N(net46));
 sg13g2_o21ai_1 \heichips25_sap3/_3585_  (.B1(\heichips25_sap3/_1161_ ),
    .Y(\heichips25_sap3/_1162_ ),
    .A1(\uio_oe_sap3[4] ),
    .A2(\heichips25_sap3/net95 ));
 sg13g2_nand4_1 \heichips25_sap3/_3586_  (.B(\heichips25_sap3/_1111_ ),
    .C(\heichips25_sap3/_1114_ ),
    .A(\heichips25_sap3/net136 ),
    .Y(\heichips25_sap3/_1163_ ),
    .D(\heichips25_sap3/_1162_ ));
 sg13g2_nor2b_1 \heichips25_sap3/_3587_  (.A(\heichips25_sap3/_1160_ ),
    .B_N(\heichips25_sap3/_1163_ ),
    .Y(\heichips25_sap3/_0108_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3588_  (.B1(\heichips25_sap3/net120 ),
    .Y(\heichips25_sap3/_1164_ ),
    .A1(\heichips25_sap3/net828 ),
    .A2(\heichips25_sap3/_1144_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3589_  (.B1(\heichips25_sap3/net136 ),
    .Y(\heichips25_sap3/_1165_ ),
    .A1(\heichips25_sap3/_1117_ ),
    .A2(\heichips25_sap3/_1164_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3590_  (.A(\heichips25_sap3/_1116_ ),
    .B(\heichips25_sap3/_1165_ ),
    .Y(\heichips25_sap3/_1166_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3591_  (.Y(\heichips25_sap3/_0109_ ),
    .B1(\heichips25_sap3/_1121_ ),
    .B2(\heichips25_sap3/_1166_ ),
    .A2(\heichips25_sap3/net100 ),
    .A1(\heichips25_sap3/_1409_ ));
 sg13g2_mux2_1 \heichips25_sap3/_3592_  (.A0(\uio_oe_sap3[6] ),
    .A1(net43),
    .S(\heichips25_sap3/_1144_ ),
    .X(\heichips25_sap3/_1167_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3593_  (.A(\heichips25_sap3/net101 ),
    .B(\heichips25_sap3/_1167_ ),
    .Y(\heichips25_sap3/_1168_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3594_  (.Y(\heichips25_sap3/_0110_ ),
    .B1(\heichips25_sap3/_1124_ ),
    .B2(\heichips25_sap3/_1168_ ),
    .A2(\heichips25_sap3/net101 ),
    .A1(\heichips25_sap3/_1417_ ));
 sg13g2_mux2_1 \heichips25_sap3/_3595_  (.A0(\uio_oe_sap3[7] ),
    .A1(net47),
    .S(\heichips25_sap3/_1144_ ),
    .X(\heichips25_sap3/_1169_ ));
 sg13g2_nor3_1 \heichips25_sap3/_3596_  (.A(\heichips25_sap3/net101 ),
    .B(\heichips25_sap3/_1131_ ),
    .C(\heichips25_sap3/_1169_ ),
    .Y(\heichips25_sap3/_1170_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3597_  (.Y(\heichips25_sap3/_0111_ ),
    .B1(\heichips25_sap3/_1130_ ),
    .B2(\heichips25_sap3/_1170_ ),
    .A2(\heichips25_sap3/net101 ),
    .A1(\heichips25_sap3/_1424_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3598_  (.A1(\heichips25_sap3/net137 ),
    .A2(\heichips25_sap3/net131 ),
    .Y(\heichips25_sap3/_1171_ ),
    .B1(\heichips25_sap3/net139 ));
 sg13g2_a21oi_1 \heichips25_sap3/_3599_  (.A1(\heichips25_sap3/net60 ),
    .A2(\heichips25_sap3/net99 ),
    .Y(\heichips25_sap3/_1172_ ),
    .B1(\heichips25_sap3/net94 ));
 sg13g2_a22oi_1 \heichips25_sap3/_3600_  (.Y(\heichips25_sap3/_1173_ ),
    .B1(\heichips25_sap3/_1172_ ),
    .B2(\heichips25_sap3/_1056_ ),
    .A2(\heichips25_sap3/net94 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][0] ));
 sg13g2_inv_1 \heichips25_sap3/_3601_  (.Y(\heichips25_sap3/_0112_ ),
    .A(\heichips25_sap3/_1173_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3602_  (.Y(\heichips25_sap3/_1174_ ),
    .A(\heichips25_sap3/_0852_ ),
    .B(\heichips25_sap3/_0888_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3603_  (.Y(\heichips25_sap3/_1175_ ),
    .A(\heichips25_sap3/_1063_ ),
    .B(\heichips25_sap3/_1174_ ));
 sg13g2_mux2_1 \heichips25_sap3/_3604_  (.A0(\heichips25_sap3/_1175_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][1] ),
    .S(\heichips25_sap3/net94 ),
    .X(\heichips25_sap3/_0113_ ));
 sg13g2_mux2_1 \heichips25_sap3/_3605_  (.A0(\heichips25_sap3/_1066_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][2] ),
    .S(\heichips25_sap3/net94 ),
    .X(\heichips25_sap3/_0114_ ));
 sg13g2_mux2_1 \heichips25_sap3/_3606_  (.A0(\heichips25_sap3/_1068_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][3] ),
    .S(\heichips25_sap3/net94 ),
    .X(\heichips25_sap3/_0115_ ));
 sg13g2_mux2_1 \heichips25_sap3/_3607_  (.A0(\heichips25_sap3/_1138_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][4] ),
    .S(\heichips25_sap3/net94 ),
    .X(\heichips25_sap3/_0116_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3608_  (.Y(\heichips25_sap3/_1176_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][5] ),
    .B(\heichips25_sap3/net94 ));
 sg13g2_o21ai_1 \heichips25_sap3/_3609_  (.B1(\heichips25_sap3/_1176_ ),
    .Y(\heichips25_sap3/_0117_ ),
    .A1(\heichips25_sap3/_1140_ ),
    .A2(\heichips25_sap3/net94 ));
 sg13g2_mux2_1 \heichips25_sap3/_3610_  (.A0(\heichips25_sap3/_1141_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][6] ),
    .S(\heichips25_sap3/_1171_ ),
    .X(\heichips25_sap3/_0118_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3611_  (.A(\heichips25_sap3/_1083_ ),
    .B(\heichips25_sap3/_1128_ ),
    .Y(\heichips25_sap3/_1177_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3612_  (.Y(\heichips25_sap3/_1178_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][7] ),
    .B(\heichips25_sap3/_1171_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3613_  (.B1(\heichips25_sap3/_1178_ ),
    .Y(\heichips25_sap3/_0119_ ),
    .A1(\heichips25_sap3/_1171_ ),
    .A2(\heichips25_sap3/_1177_ ));
 sg13g2_nand3_1 \heichips25_sap3/_3614_  (.B(\heichips25_sap3/_0876_ ),
    .C(\heichips25_sap3/_1056_ ),
    .A(\heichips25_sap3/net140 ),
    .Y(\heichips25_sap3/_1179_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3615_  (.B1(\heichips25_sap3/_1179_ ),
    .Y(\heichips25_sap3/_0120_ ),
    .A1(\heichips25_sap3/_1394_ ),
    .A2(\heichips25_sap3/net141 ));
 sg13g2_nor3_1 \heichips25_sap3/_3616_  (.A(\heichips25_sap3/net102 ),
    .B(\heichips25_sap3/_1061_ ),
    .C(\heichips25_sap3/_1093_ ),
    .Y(\heichips25_sap3/_1180_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3617_  (.A1(\heichips25_sap3/_1388_ ),
    .A2(\heichips25_sap3/net102 ),
    .Y(\heichips25_sap3/_0121_ ),
    .B1(\heichips25_sap3/_1180_ ));
 sg13g2_and2_1 \heichips25_sap3/_3618_  (.A(\heichips25_sap3/net141 ),
    .B(\heichips25_sap3/_1064_ ),
    .X(\heichips25_sap3/_1181_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3619_  (.Y(\heichips25_sap3/_0122_ ),
    .B1(\heichips25_sap3/_0929_ ),
    .B2(\heichips25_sap3/_1181_ ),
    .A2(\heichips25_sap3/net102 ),
    .A1(\heichips25_sap3/_1378_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3620_  (.A(\heichips25_sap3/net102 ),
    .B(\heichips25_sap3/_1067_ ),
    .Y(\heichips25_sap3/_1182_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3621_  (.Y(\heichips25_sap3/_0123_ ),
    .B1(\heichips25_sap3/_1106_ ),
    .B2(\heichips25_sap3/_1182_ ),
    .A2(\heichips25_sap3/net102 ),
    .A1(\heichips25_sap3/_1371_ ));
 sg13g2_nor3_1 \heichips25_sap3/_3622_  (.A(\heichips25_sap3/net102 ),
    .B(\heichips25_sap3/_0984_ ),
    .C(\heichips25_sap3/_1069_ ),
    .Y(\heichips25_sap3/_1183_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3623_  (.Y(\heichips25_sap3/_0124_ ),
    .B1(\heichips25_sap3/_1111_ ),
    .B2(\heichips25_sap3/_1183_ ),
    .A2(\heichips25_sap3/net102 ),
    .A1(\heichips25_sap3/_1403_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3624_  (.A(\heichips25_sap3/net102 ),
    .B(\heichips25_sap3/_1073_ ),
    .Y(\heichips25_sap3/_1184_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3625_  (.Y(\heichips25_sap3/_0125_ ),
    .B1(\heichips25_sap3/_1121_ ),
    .B2(\heichips25_sap3/_1184_ ),
    .A2(\heichips25_sap3/net103 ),
    .A1(\heichips25_sap3/_1408_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3626_  (.A(\heichips25_sap3/net103 ),
    .B(\heichips25_sap3/_1078_ ),
    .Y(\heichips25_sap3/_1185_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3627_  (.Y(\heichips25_sap3/_0126_ ),
    .B1(\heichips25_sap3/_1122_ ),
    .B2(\heichips25_sap3/_1185_ ),
    .A2(\heichips25_sap3/net103 ),
    .A1(\heichips25_sap3/_1416_ ));
 sg13g2_and2_1 \heichips25_sap3/_3628_  (.A(\heichips25_sap3/net142 ),
    .B(\heichips25_sap3/_1082_ ),
    .X(\heichips25_sap3/_1186_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3629_  (.Y(\heichips25_sap3/_0127_ ),
    .B1(\heichips25_sap3/_1130_ ),
    .B2(\heichips25_sap3/_1186_ ),
    .A2(\heichips25_sap3/net103 ),
    .A1(\heichips25_sap3/_1423_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3630_  (.A1(\heichips25_sap3/net142 ),
    .A2(\heichips25_sap3/_0881_ ),
    .Y(\heichips25_sap3/_1187_ ),
    .B1(\heichips25_sap3/net132 ));
 sg13g2_a21oi_1 \heichips25_sap3/_3631_  (.A1(\heichips25_sap3/net60 ),
    .A2(\heichips25_sap3/net99 ),
    .Y(\heichips25_sap3/_1188_ ),
    .B1(\heichips25_sap3/net93 ));
 sg13g2_a22oi_1 \heichips25_sap3/_3632_  (.Y(\heichips25_sap3/_1189_ ),
    .B1(\heichips25_sap3/_1188_ ),
    .B2(\heichips25_sap3/_1056_ ),
    .A2(\heichips25_sap3/net93 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][0] ));
 sg13g2_inv_1 \heichips25_sap3/_3633_  (.Y(\heichips25_sap3/_0128_ ),
    .A(\heichips25_sap3/_1189_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3634_  (.Y(\heichips25_sap3/_1190_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][1] ),
    .B(\heichips25_sap3/net93 ));
 sg13g2_o21ai_1 \heichips25_sap3/_3635_  (.B1(\heichips25_sap3/_1190_ ),
    .Y(\heichips25_sap3/_0129_ ),
    .A1(\heichips25_sap3/_1063_ ),
    .A2(\heichips25_sap3/net93 ));
 sg13g2_mux2_1 \heichips25_sap3/_3636_  (.A0(\heichips25_sap3/_1066_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][2] ),
    .S(\heichips25_sap3/net93 ),
    .X(\heichips25_sap3/_0130_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3637_  (.A1(\heichips25_sap3/_0888_ ),
    .A2(\heichips25_sap3/_1159_ ),
    .Y(\heichips25_sap3/_1191_ ),
    .B1(\heichips25_sap3/_1068_ ));
 sg13g2_mux2_1 \heichips25_sap3/_3638_  (.A0(\heichips25_sap3/_1068_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][3] ),
    .S(\heichips25_sap3/net93 ),
    .X(\heichips25_sap3/_0131_ ));
 sg13g2_mux2_1 \heichips25_sap3/_3639_  (.A0(\heichips25_sap3/_1138_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][4] ),
    .S(\heichips25_sap3/net93 ),
    .X(\heichips25_sap3/_0132_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3640_  (.Y(\heichips25_sap3/_1192_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][5] ),
    .B(\heichips25_sap3/net93 ));
 sg13g2_o21ai_1 \heichips25_sap3/_3641_  (.B1(\heichips25_sap3/_1192_ ),
    .Y(\heichips25_sap3/_0133_ ),
    .A1(\heichips25_sap3/_1140_ ),
    .A2(\heichips25_sap3/_1187_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3642_  (.A1(\heichips25_sap3/_0794_ ),
    .A2(\heichips25_sap3/_0868_ ),
    .Y(\heichips25_sap3/_1193_ ),
    .B1(\heichips25_sap3/_0889_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3643_  (.A1(\heichips25_sap3/_0869_ ),
    .A2(\heichips25_sap3/_1193_ ),
    .Y(\heichips25_sap3/_1194_ ),
    .B1(\heichips25_sap3/_1078_ ));
 sg13g2_mux2_1 \heichips25_sap3/_3644_  (.A0(\heichips25_sap3/_1141_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][6] ),
    .S(\heichips25_sap3/_1187_ ),
    .X(\heichips25_sap3/_0134_ ));
 sg13g2_mux2_1 \heichips25_sap3/_3645_  (.A0(\heichips25_sap3/_1083_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][7] ),
    .S(\heichips25_sap3/_1187_ ),
    .X(\heichips25_sap3/_0135_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3646_  (.A(\heichips25_sap3/net49 ),
    .B(\heichips25_sap3/_0889_ ),
    .Y(\heichips25_sap3/_1195_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3647_  (.B1(\heichips25_sap3/_1195_ ),
    .Y(\heichips25_sap3/_1196_ ),
    .A1(\heichips25_sap3/_0777_ ),
    .A2(\heichips25_sap3/_0870_ ));
 sg13g2_nor3_1 \heichips25_sap3/_3648_  (.A(\uio_oe_sap3[0] ),
    .B(\heichips25_sap3/net98 ),
    .C(\heichips25_sap3/_1053_ ),
    .Y(\heichips25_sap3/_1197_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_3649_  (.B2(\heichips25_sap3/_1197_ ),
    .C1(\heichips25_sap3/net112 ),
    .B1(\heichips25_sap3/_1196_ ),
    .A1(\heichips25_sap3/net98 ),
    .Y(\heichips25_sap3/_1198_ ),
    .A2(\heichips25_sap3/_0875_ ));
 sg13g2_a21o_1 \heichips25_sap3/_3650_  (.A2(\heichips25_sap3/net112 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][0] ),
    .B1(\heichips25_sap3/_1198_ ),
    .X(\heichips25_sap3/_0136_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3651_  (.A1(\heichips25_sap3/net48 ),
    .A2(\heichips25_sap3/net51 ),
    .Y(\heichips25_sap3/_1199_ ),
    .B1(\heichips25_sap3/_0889_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3652_  (.B1(\heichips25_sap3/_1199_ ),
    .Y(\heichips25_sap3/_1200_ ),
    .A1(\heichips25_sap3/net48 ),
    .A2(\heichips25_sap3/net51 ));
 sg13g2_and3_1 \heichips25_sap3/_3653_  (.X(\heichips25_sap3/_1201_ ),
    .A(\heichips25_sap3/_0327_ ),
    .B(\heichips25_sap3/net146 ),
    .C(\heichips25_sap3/_1200_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3654_  (.Y(\heichips25_sap3/_0137_ ),
    .B1(\heichips25_sap3/_1095_ ),
    .B2(\heichips25_sap3/_1201_ ),
    .A2(\heichips25_sap3/net112 ),
    .A1(\heichips25_sap3/_1387_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3655_  (.A1(\heichips25_sap3/net48 ),
    .A2(\heichips25_sap3/net51 ),
    .Y(\heichips25_sap3/_1202_ ),
    .B1(\heichips25_sap3/net50 ));
 sg13g2_nor2_1 \heichips25_sap3/_3656_  (.A(\heichips25_sap3/_0889_ ),
    .B(\heichips25_sap3/_1202_ ),
    .Y(\heichips25_sap3/_1203_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_3657_  (.Y(\heichips25_sap3/_1204_ ),
    .B(\heichips25_sap3/net119 ),
    .A_N(\uio_oe_sap3[2] ));
 sg13g2_a221oi_1 \heichips25_sap3/_3658_  (.B2(\heichips25_sap3/_1104_ ),
    .C1(\heichips25_sap3/net112 ),
    .B1(\heichips25_sap3/_1204_ ),
    .A1(\heichips25_sap3/_0927_ ),
    .Y(\heichips25_sap3/_1205_ ),
    .A2(\heichips25_sap3/_1203_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3659_  (.Y(\heichips25_sap3/_0138_ ),
    .B1(\heichips25_sap3/_0929_ ),
    .B2(\heichips25_sap3/_1205_ ),
    .A2(\heichips25_sap3/net112 ),
    .A1(\heichips25_sap3/_1377_ ));
 sg13g2_xor2_1 \heichips25_sap3/_3660_  (.B(\heichips25_sap3/_0943_ ),
    .A(\heichips25_sap3/_0927_ ),
    .X(\heichips25_sap3/_1206_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3661_  (.A1(\heichips25_sap3/net146 ),
    .A2(\heichips25_sap3/_1206_ ),
    .Y(\heichips25_sap3/_1207_ ),
    .B1(\heichips25_sap3/_0889_ ));
 sg13g2_nor3_1 \heichips25_sap3/_3662_  (.A(\uio_oe_sap3[3] ),
    .B(\heichips25_sap3/net112 ),
    .C(\heichips25_sap3/_1207_ ),
    .Y(\heichips25_sap3/_1208_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3663_  (.Y(\heichips25_sap3/_0139_ ),
    .B1(\heichips25_sap3/_1106_ ),
    .B2(\heichips25_sap3/_1208_ ),
    .A2(\heichips25_sap3/net112 ),
    .A1(\heichips25_sap3/_1370_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3664_  (.B1(\heichips25_sap3/net146 ),
    .Y(\heichips25_sap3/_1209_ ),
    .A1(\uio_oe_sap3[4] ),
    .A2(\heichips25_sap3/_0732_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3665_  (.B1(\heichips25_sap3/_0969_ ),
    .Y(\heichips25_sap3/_1210_ ),
    .A1(\heichips25_sap3/_0945_ ),
    .A2(\heichips25_sap3/_0965_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_3666_  (.B2(\heichips25_sap3/_0888_ ),
    .C1(\heichips25_sap3/_1209_ ),
    .B1(\heichips25_sap3/_1210_ ),
    .A1(\heichips25_sap3/net96 ),
    .Y(\heichips25_sap3/_1211_ ),
    .A2(\heichips25_sap3/_0971_ ));
 sg13g2_a21o_1 \heichips25_sap3/_3667_  (.A2(\heichips25_sap3/net111 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][4] ),
    .B1(\heichips25_sap3/_1211_ ),
    .X(\heichips25_sap3/_0140_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3668_  (.A(\heichips25_sap3/net828 ),
    .B(\heichips25_sap3/net111 ),
    .Y(\heichips25_sap3/_1212_ ));
 sg13g2_xnor2_1 \heichips25_sap3/_3669_  (.Y(\heichips25_sap3/_1213_ ),
    .A(\heichips25_sap3/_0969_ ),
    .B(\heichips25_sap3/_0991_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3670_  (.B1(\heichips25_sap3/_0888_ ),
    .Y(\heichips25_sap3/_1214_ ),
    .A1(\heichips25_sap3/net111 ),
    .A2(\heichips25_sap3/_1213_ ));
 sg13g2_and2_1 \heichips25_sap3/_3671_  (.A(\heichips25_sap3/_1212_ ),
    .B(\heichips25_sap3/_1214_ ),
    .X(\heichips25_sap3/_1215_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3672_  (.Y(\heichips25_sap3/_0141_ ),
    .B1(\heichips25_sap3/_1121_ ),
    .B2(\heichips25_sap3/_1215_ ),
    .A2(\heichips25_sap3/net111 ),
    .A1(\heichips25_sap3/_1407_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3673_  (.Y(\heichips25_sap3/_1216_ ),
    .A(\heichips25_sap3/_0992_ ),
    .B(\heichips25_sap3/_1015_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3674_  (.A(\heichips25_sap3/_0889_ ),
    .B(\heichips25_sap3/_1017_ ),
    .Y(\heichips25_sap3/_1217_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_3675_  (.Y(\heichips25_sap3/_1218_ ),
    .B(\heichips25_sap3/net146 ),
    .A_N(\uio_oe_sap3[6] ));
 sg13g2_a21oi_1 \heichips25_sap3/_3676_  (.A1(\heichips25_sap3/_1216_ ),
    .A2(\heichips25_sap3/_1217_ ),
    .Y(\heichips25_sap3/_1219_ ),
    .B1(\heichips25_sap3/_1218_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3677_  (.Y(\heichips25_sap3/_0142_ ),
    .B1(\heichips25_sap3/_1122_ ),
    .B2(\heichips25_sap3/_1219_ ),
    .A2(\heichips25_sap3/net111 ),
    .A1(\heichips25_sap3/_1415_ ));
 sg13g2_xor2_1 \heichips25_sap3/_3678_  (.B(\heichips25_sap3/_1036_ ),
    .A(\heichips25_sap3/_1017_ ),
    .X(\heichips25_sap3/_1220_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_3679_  (.Y(\heichips25_sap3/_1221_ ),
    .B(\heichips25_sap3/net149 ),
    .A_N(\uio_oe_sap3[7] ));
 sg13g2_a21oi_1 \heichips25_sap3/_3680_  (.A1(\heichips25_sap3/_0888_ ),
    .A2(\heichips25_sap3/_1220_ ),
    .Y(\heichips25_sap3/_1222_ ),
    .B1(\heichips25_sap3/_1221_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3681_  (.Y(\heichips25_sap3/_0143_ ),
    .B1(\heichips25_sap3/_1129_ ),
    .B2(\heichips25_sap3/_1222_ ),
    .A2(\heichips25_sap3/net111 ),
    .A1(\heichips25_sap3/_1422_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3682_  (.A1(\heichips25_sap3/net60 ),
    .A2(\heichips25_sap3/net99 ),
    .Y(\heichips25_sap3/_1223_ ),
    .B1(\heichips25_sap3/net113 ));
 sg13g2_a22oi_1 \heichips25_sap3/_3683_  (.Y(\heichips25_sap3/_1224_ ),
    .B1(\heichips25_sap3/_1056_ ),
    .B2(\heichips25_sap3/_1223_ ),
    .A2(\heichips25_sap3/net113 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][0] ));
 sg13g2_inv_1 \heichips25_sap3/_3684_  (.Y(\heichips25_sap3/_0144_ ),
    .A(\heichips25_sap3/_1224_ ));
 sg13g2_mux2_1 \heichips25_sap3/_3685_  (.A0(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][1] ),
    .A1(\heichips25_sap3/_1175_ ),
    .S(\heichips25_sap3/net147 ),
    .X(\heichips25_sap3/_0145_ ));
 sg13g2_mux2_1 \heichips25_sap3/_3686_  (.A0(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][2] ),
    .A1(\heichips25_sap3/_1066_ ),
    .S(\heichips25_sap3/net147 ),
    .X(\heichips25_sap3/_0146_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3687_  (.Y(\heichips25_sap3/_1225_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][3] ),
    .B(\heichips25_sap3/net113 ));
 sg13g2_o21ai_1 \heichips25_sap3/_3688_  (.B1(\heichips25_sap3/_1225_ ),
    .Y(\heichips25_sap3/_0147_ ),
    .A1(\heichips25_sap3/net112 ),
    .A2(\heichips25_sap3/_1191_ ));
 sg13g2_nor4_1 \heichips25_sap3/_3689_  (.A(\heichips25_sap3/net111 ),
    .B(\heichips25_sap3/_0984_ ),
    .C(\heichips25_sap3/_1069_ ),
    .D(\heichips25_sap3/_1137_ ),
    .Y(\heichips25_sap3/_1226_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3690_  (.A1(\heichips25_sap3/_1402_ ),
    .A2(\heichips25_sap3/net113 ),
    .Y(\heichips25_sap3/_0148_ ),
    .B1(\heichips25_sap3/_1226_ ));
 sg13g2_xnor2_1 \heichips25_sap3/_3691_  (.Y(\heichips25_sap3/_1227_ ),
    .A(\heichips25_sap3/_0802_ ),
    .B(\heichips25_sap3/_0867_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3692_  (.A1(\heichips25_sap3/_0888_ ),
    .A2(\heichips25_sap3/_1227_ ),
    .Y(\heichips25_sap3/_1228_ ),
    .B1(\heichips25_sap3/net113 ));
 sg13g2_a22oi_1 \heichips25_sap3/_3693_  (.Y(\heichips25_sap3/_0149_ ),
    .B1(\heichips25_sap3/_1140_ ),
    .B2(\heichips25_sap3/_1228_ ),
    .A2(\heichips25_sap3/_0755_ ),
    .A1(\heichips25_sap3/_1406_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3694_  (.A(\heichips25_sap3/net111 ),
    .B(\heichips25_sap3/_1079_ ),
    .Y(\heichips25_sap3/_1229_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3695_  (.Y(\heichips25_sap3/_0150_ ),
    .B1(\heichips25_sap3/_1194_ ),
    .B2(\heichips25_sap3/_1229_ ),
    .A2(\heichips25_sap3/net113 ),
    .A1(\heichips25_sap3/_1414_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3696_  (.Y(\heichips25_sap3/_1230_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][7] ),
    .B(\heichips25_sap3/_0755_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3697_  (.B1(\heichips25_sap3/_1230_ ),
    .Y(\heichips25_sap3/_0151_ ),
    .A1(\heichips25_sap3/_0755_ ),
    .A2(\heichips25_sap3/_1177_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3698_  (.Y(\heichips25_sap3/_1231_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][0] ),
    .B(\heichips25_sap3/net115 ));
 sg13g2_nand2_1 \heichips25_sap3/_3699_  (.Y(\heichips25_sap3/_1232_ ),
    .A(\heichips25_sap3/net116 ),
    .B(\heichips25_sap3/_0876_ ));
 sg13g2_nor3_1 \heichips25_sap3/_3700_  (.A(\uio_oe_sap3[0] ),
    .B(\heichips25_sap3/_1055_ ),
    .C(\heichips25_sap3/_1086_ ),
    .Y(\heichips25_sap3/_1233_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3701_  (.B1(\heichips25_sap3/_1231_ ),
    .Y(\heichips25_sap3/_0152_ ),
    .A1(\heichips25_sap3/_1232_ ),
    .A2(\heichips25_sap3/_1233_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3702_  (.A(\uio_oe_sap3[1] ),
    .B(\heichips25_sap3/net115 ),
    .Y(\heichips25_sap3/_1234_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3703_  (.Y(\heichips25_sap3/_0153_ ),
    .B1(\heichips25_sap3/_1095_ ),
    .B2(\heichips25_sap3/_1234_ ),
    .A2(\heichips25_sap3/net115 ),
    .A1(\heichips25_sap3/_1386_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3704_  (.A1(\heichips25_sap3/_1100_ ),
    .A2(\heichips25_sap3/_1204_ ),
    .Y(\heichips25_sap3/_1235_ ),
    .B1(\heichips25_sap3/net115 ));
 sg13g2_a22oi_1 \heichips25_sap3/_3705_  (.Y(\heichips25_sap3/_0154_ ),
    .B1(\heichips25_sap3/_0929_ ),
    .B2(\heichips25_sap3/_1235_ ),
    .A2(\heichips25_sap3/net115 ),
    .A1(\heichips25_sap3/_1376_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3706_  (.A(\uio_oe_sap3[3] ),
    .B(\heichips25_sap3/net115 ),
    .Y(\heichips25_sap3/_1236_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3707_  (.Y(\heichips25_sap3/_0155_ ),
    .B1(\heichips25_sap3/_1107_ ),
    .B2(\heichips25_sap3/_1236_ ),
    .A2(\heichips25_sap3/net115 ),
    .A1(\heichips25_sap3/_1369_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3708_  (.A(\uio_oe_sap3[4] ),
    .B(\heichips25_sap3/net114 ),
    .Y(\heichips25_sap3/_1237_ ));
 sg13g2_and2_1 \heichips25_sap3/_3709_  (.A(\heichips25_sap3/_1114_ ),
    .B(\heichips25_sap3/_1237_ ),
    .X(\heichips25_sap3/_1238_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3710_  (.Y(\heichips25_sap3/_0156_ ),
    .B1(\heichips25_sap3/_1111_ ),
    .B2(\heichips25_sap3/_1238_ ),
    .A2(\heichips25_sap3/net114 ),
    .A1(\heichips25_sap3/_1401_ ));
 sg13g2_nor3_1 \heichips25_sap3/_3711_  (.A(\heichips25_sap3/net828 ),
    .B(\heichips25_sap3/net114 ),
    .C(\heichips25_sap3/_1116_ ),
    .Y(\heichips25_sap3/_1239_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3712_  (.Y(\heichips25_sap3/_0157_ ),
    .B1(\heichips25_sap3/_1121_ ),
    .B2(\heichips25_sap3/_1239_ ),
    .A2(\heichips25_sap3/net114 ),
    .A1(\heichips25_sap3/_1405_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3713_  (.A(\uio_oe_sap3[6] ),
    .B(\heichips25_sap3/net114 ),
    .Y(\heichips25_sap3/_1240_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3714_  (.Y(\heichips25_sap3/_0158_ ),
    .B1(\heichips25_sap3/_1124_ ),
    .B2(\heichips25_sap3/_1240_ ),
    .A2(\heichips25_sap3/net114 ),
    .A1(\heichips25_sap3/_1413_ ));
 sg13g2_nor3_1 \heichips25_sap3/_3715_  (.A(\uio_oe_sap3[7] ),
    .B(\heichips25_sap3/net114 ),
    .C(\heichips25_sap3/_1131_ ),
    .Y(\heichips25_sap3/_1241_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3716_  (.Y(\heichips25_sap3/_0159_ ),
    .B1(\heichips25_sap3/_1129_ ),
    .B2(\heichips25_sap3/_1241_ ),
    .A2(\heichips25_sap3/net114 ),
    .A1(\heichips25_sap3/_1421_ ));
 sg13g2_nand3_1 \heichips25_sap3/_3717_  (.B(\heichips25_sap3/_1056_ ),
    .C(\heichips25_sap3/_1057_ ),
    .A(\heichips25_sap3/net117 ),
    .Y(\heichips25_sap3/_1242_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3718_  (.B1(\heichips25_sap3/_1242_ ),
    .Y(\heichips25_sap3/_0160_ ),
    .A1(\heichips25_sap3/_1393_ ),
    .A2(\heichips25_sap3/net117 ));
 sg13g2_mux2_1 \heichips25_sap3/_3719_  (.A0(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][1] ),
    .A1(\heichips25_sap3/_1175_ ),
    .S(\heichips25_sap3/net117 ),
    .X(\heichips25_sap3/_0161_ ));
 sg13g2_mux2_1 \heichips25_sap3/_3720_  (.A0(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][2] ),
    .A1(\heichips25_sap3/_1066_ ),
    .S(\heichips25_sap3/net117 ),
    .X(\heichips25_sap3/_0162_ ));
 sg13g2_mux2_1 \heichips25_sap3/_3721_  (.A0(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][3] ),
    .A1(\heichips25_sap3/_1068_ ),
    .S(\heichips25_sap3/net117 ),
    .X(\heichips25_sap3/_0163_ ));
 sg13g2_mux2_1 \heichips25_sap3/_3722_  (.A0(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][4] ),
    .A1(\heichips25_sap3/_1138_ ),
    .S(\heichips25_sap3/net117 ),
    .X(\heichips25_sap3/_0164_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3723_  (.Y(\heichips25_sap3/_1243_ ),
    .A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][5] ),
    .B(\heichips25_sap3/_0753_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3724_  (.B1(\heichips25_sap3/_1243_ ),
    .Y(\heichips25_sap3/_0165_ ),
    .A1(\heichips25_sap3/_0753_ ),
    .A2(\heichips25_sap3/_1140_ ));
 sg13g2_mux2_1 \heichips25_sap3/_3725_  (.A0(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][6] ),
    .A1(\heichips25_sap3/_1141_ ),
    .S(\heichips25_sap3/net118 ),
    .X(\heichips25_sap3/_0166_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3726_  (.A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][7] ),
    .B(\heichips25_sap3/net118 ),
    .Y(\heichips25_sap3/_1244_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3727_  (.A1(\heichips25_sap3/net118 ),
    .A2(\heichips25_sap3/_1177_ ),
    .Y(\heichips25_sap3/_0167_ ),
    .B1(\heichips25_sap3/_1244_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3728_  (.Y(\heichips25_sap3/_1245_ ),
    .A(\heichips25_sap3/_1360_ ),
    .B(\heichips25_sap3/net832 ));
 sg13g2_nand2_1 \heichips25_sap3/_3729_  (.Y(\heichips25_sap3/_1246_ ),
    .A(\heichips25_sap3/_0291_ ),
    .B(\heichips25_sap3/_1245_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3730_  (.A(\heichips25_sap3/net1058 ),
    .B(\heichips25_sap3/_1246_ ),
    .Y(\heichips25_sap3/_1247_ ));
 sg13g2_nand3b_1 \heichips25_sap3/_3731_  (.B(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos[1] ),
    .C(\heichips25_sap3/net1031 ),
    .Y(\heichips25_sap3/_1248_ ),
    .A_N(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos[0] ));
 sg13g2_a21oi_1 \heichips25_sap3/_3732_  (.A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos[0] ),
    .A2(\heichips25_sap3/_1426_ ),
    .Y(\heichips25_sap3/_1249_ ),
    .B1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos[1] ));
 sg13g2_o21ai_1 \heichips25_sap3/_3733_  (.B1(\heichips25_sap3/_1249_ ),
    .Y(\heichips25_sap3/_1250_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos[0] ),
    .A2(\heichips25_sap3/net1011 ));
 sg13g2_a21oi_1 \heichips25_sap3/_3734_  (.A1(\heichips25_sap3/_1248_ ),
    .A2(\heichips25_sap3/_1250_ ),
    .Y(\heichips25_sap3/_1251_ ),
    .B1(\heichips25_sap3/_1432_ ));
 sg13g2_mux4_1 \heichips25_sap3/_3735_  (.S0(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos[0] ),
    .A0(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[1] ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[2] ),
    .A2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[3] ),
    .A3(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[4] ),
    .S1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos[1] ),
    .X(\heichips25_sap3/_1252_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_3736_  (.B2(\heichips25_sap3/_1252_ ),
    .C1(\heichips25_sap3/_1251_ ),
    .B1(\heichips25_sap3/_0290_ ),
    .A1(\heichips25_sap3/_1360_ ),
    .Y(\heichips25_sap3/_1253_ ),
    .A2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[0] ));
 sg13g2_a21oi_1 \heichips25_sap3/_3737_  (.A1(\heichips25_sap3/_1246_ ),
    .A2(\heichips25_sap3/_1253_ ),
    .Y(\heichips25_sap3/_0168_ ),
    .B1(\heichips25_sap3/_1247_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3738_  (.A1(\heichips25_sap3/_1429_ ),
    .A2(\heichips25_sap3/net339 ),
    .Y(\heichips25_sap3/_0169_ ),
    .B1(\heichips25_sap3/net832 ));
 sg13g2_nor2_1 \heichips25_sap3/_3739_  (.A(\heichips25_sap3/net1130 ),
    .B(\heichips25_sap3/net1176 ),
    .Y(\heichips25_sap3/_1254_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3740_  (.A1(\heichips25_sap3/net1176 ),
    .A2(\heichips25_sap3/_1246_ ),
    .Y(\heichips25_sap3/_0170_ ),
    .B1(\heichips25_sap3/_1254_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3741_  (.A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos[0] ),
    .A2(\heichips25_sap3/_1246_ ),
    .Y(\heichips25_sap3/_1255_ ),
    .B1(\heichips25_sap3/net1162 ));
 sg13g2_a21oi_1 \heichips25_sap3/_3742_  (.A1(\heichips25_sap3/_0289_ ),
    .A2(\heichips25_sap3/_1246_ ),
    .Y(\heichips25_sap3/_0171_ ),
    .B1(\heichips25_sap3/net1163 ));
 sg13g2_nand2_1 \heichips25_sap3/_3743_  (.Y(\heichips25_sap3/_1256_ ),
    .A(\heichips25_sap3/net835 ),
    .B(\heichips25_sap3/_1245_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3744_  (.B1(\heichips25_sap3/net836 ),
    .Y(\heichips25_sap3/_0172_ ),
    .A1(\heichips25_sap3/_1360_ ),
    .A2(\heichips25_sap3/_1431_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_3745_  (.Y(\heichips25_sap3/_1257_ ),
    .B(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.word_index[2] ),
    .A_N(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.word_index[3] ));
 sg13g2_nand2_1 \heichips25_sap3/_3746_  (.Y(\heichips25_sap3/_1258_ ),
    .A(\heichips25_sap3/_1428_ ),
    .B(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.word_index[1] ));
 sg13g2_nor2_1 \heichips25_sap3/_3747_  (.A(\heichips25_sap3/_1257_ ),
    .B(\heichips25_sap3/_1258_ ),
    .Y(\heichips25_sap3/_1259_ ));
 sg13g2_nand2_1 \heichips25_sap3/_3748_  (.Y(\heichips25_sap3/_1260_ ),
    .A(\heichips25_sap3/net1197 ),
    .B(\heichips25_sap3/net1178 ));
 sg13g2_nor2_1 \heichips25_sap3/_3749_  (.A(\heichips25_sap3/_1257_ ),
    .B(\heichips25_sap3/_1260_ ),
    .Y(\heichips25_sap3/_1261_ ));
 sg13g2_inv_1 \heichips25_sap3/_3750_  (.Y(\heichips25_sap3/_1262_ ),
    .A(\heichips25_sap3/net293 ));
 sg13g2_a22oi_1 \heichips25_sap3/_3751_  (.Y(\heichips25_sap3/_1263_ ),
    .B1(\heichips25_sap3/net293 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][0] ),
    .A2(\heichips25_sap3/_1259_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][0] ));
 sg13g2_nand2b_1 \heichips25_sap3/_3752_  (.Y(\heichips25_sap3/_1264_ ),
    .B(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.word_index[3] ),
    .A_N(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.word_index[2] ));
 sg13g2_nor3_1 \heichips25_sap3/_3753_  (.A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.word_index[0] ),
    .B(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.word_index[1] ),
    .C(\heichips25_sap3/_1264_ ),
    .Y(\heichips25_sap3/_1265_ ));
 sg13g2_nor3_1 \heichips25_sap3/_3754_  (.A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.word_index[3] ),
    .B(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.word_index[2] ),
    .C(\heichips25_sap3/_1260_ ),
    .Y(\heichips25_sap3/_1266_ ));
 sg13g2_inv_1 \heichips25_sap3/_3755_  (.Y(\heichips25_sap3/_1267_ ),
    .A(\heichips25_sap3/net292 ));
 sg13g2_a22oi_1 \heichips25_sap3/_3756_  (.Y(\heichips25_sap3/_1268_ ),
    .B1(\heichips25_sap3/net292 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][0] ),
    .A2(\heichips25_sap3/_1265_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][0] ));
 sg13g2_nand2_1 \heichips25_sap3/_3757_  (.Y(\heichips25_sap3/_1269_ ),
    .A(\heichips25_sap3/_1263_ ),
    .B(\heichips25_sap3/_1268_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3758_  (.A(\heichips25_sap3/_1260_ ),
    .B(\heichips25_sap3/_1264_ ),
    .Y(\heichips25_sap3/_1270_ ));
 sg13g2_nand2b_1 \heichips25_sap3/_3759_  (.Y(\heichips25_sap3/_1271_ ),
    .B(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.word_index[0] ),
    .A_N(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.word_index[1] ));
 sg13g2_nor2_1 \heichips25_sap3/_3760_  (.A(\heichips25_sap3/_1257_ ),
    .B(\heichips25_sap3/_1271_ ),
    .Y(\heichips25_sap3/_1272_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3761_  (.Y(\heichips25_sap3/_1273_ ),
    .B1(\heichips25_sap3/_1272_ ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][0] ),
    .A2(\heichips25_sap3/_1270_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][0] ));
 sg13g2_nor3_1 \heichips25_sap3/_3762_  (.A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.word_index[3] ),
    .B(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.word_index[2] ),
    .C(\heichips25_sap3/_1271_ ),
    .Y(\heichips25_sap3/_1274_ ));
 sg13g2_nor4_1 \heichips25_sap3/_3763_  (.A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.word_index[0] ),
    .B(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.word_index[1] ),
    .C(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.word_index[3] ),
    .D(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.word_index[2] ),
    .Y(\heichips25_sap3/_1275_ ));
 sg13g2_a21o_1 \heichips25_sap3/_3764_  (.A2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.word_index[2] ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.word_index[3] ),
    .B1(\heichips25_sap3/_1275_ ),
    .X(\heichips25_sap3/_1276_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3765_  (.A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][0] ),
    .A2(\heichips25_sap3/_1274_ ),
    .Y(\heichips25_sap3/_1277_ ),
    .B1(\heichips25_sap3/net290 ));
 sg13g2_nor2_1 \heichips25_sap3/_3766_  (.A(\heichips25_sap3/_1264_ ),
    .B(\heichips25_sap3/_1271_ ),
    .Y(\heichips25_sap3/_1278_ ));
 sg13g2_nor3_1 \heichips25_sap3/_3767_  (.A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.word_index[0] ),
    .B(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.word_index[1] ),
    .C(\heichips25_sap3/_1257_ ),
    .Y(\heichips25_sap3/_1279_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3768_  (.Y(\heichips25_sap3/_1280_ ),
    .B1(\heichips25_sap3/_1279_ ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][0] ),
    .A2(\heichips25_sap3/_1278_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][0] ));
 sg13g2_nor2_1 \heichips25_sap3/_3769_  (.A(\heichips25_sap3/_1258_ ),
    .B(\heichips25_sap3/_1264_ ),
    .Y(\heichips25_sap3/_1281_ ));
 sg13g2_nor3_1 \heichips25_sap3/_3770_  (.A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.word_index[3] ),
    .B(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.word_index[2] ),
    .C(\heichips25_sap3/_1258_ ),
    .Y(\heichips25_sap3/_1282_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3771_  (.Y(\heichips25_sap3/_1283_ ),
    .B1(\heichips25_sap3/_1282_ ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][0] ),
    .A2(\heichips25_sap3/_1281_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][0] ));
 sg13g2_nand4_1 \heichips25_sap3/_3772_  (.B(\heichips25_sap3/_1277_ ),
    .C(\heichips25_sap3/_1280_ ),
    .A(\heichips25_sap3/_1273_ ),
    .Y(\heichips25_sap3/_1284_ ),
    .D(\heichips25_sap3/_1283_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3773_  (.A1(\heichips25_sap3/_1392_ ),
    .A2(\heichips25_sap3/net290 ),
    .Y(\heichips25_sap3/_1285_ ),
    .B1(\heichips25_sap3/net339 ));
 sg13g2_o21ai_1 \heichips25_sap3/_3774_  (.B1(\heichips25_sap3/_1285_ ),
    .Y(\heichips25_sap3/_1286_ ),
    .A1(\heichips25_sap3/_1269_ ),
    .A2(\heichips25_sap3/_1284_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3775_  (.B1(\heichips25_sap3/_1286_ ),
    .Y(\heichips25_sap3/_0173_ ),
    .A1(\heichips25_sap3/_1427_ ),
    .A2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.state[0] ));
 sg13g2_a22oi_1 \heichips25_sap3/_3776_  (.Y(\heichips25_sap3/_1287_ ),
    .B1(\heichips25_sap3/_1278_ ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][1] ),
    .A2(\heichips25_sap3/_1259_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][1] ));
 sg13g2_a22oi_1 \heichips25_sap3/_3777_  (.Y(\heichips25_sap3/_1288_ ),
    .B1(\heichips25_sap3/_1282_ ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][1] ),
    .A2(\heichips25_sap3/_1265_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][1] ));
 sg13g2_a21oi_1 \heichips25_sap3/_3778_  (.A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][1] ),
    .A2(\heichips25_sap3/_1279_ ),
    .Y(\heichips25_sap3/_1289_ ),
    .B1(\heichips25_sap3/net290 ));
 sg13g2_a22oi_1 \heichips25_sap3/_3779_  (.Y(\heichips25_sap3/_1290_ ),
    .B1(\heichips25_sap3/net292 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][1] ),
    .A2(\heichips25_sap3/net293 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][1] ));
 sg13g2_a22oi_1 \heichips25_sap3/_3780_  (.Y(\heichips25_sap3/_1291_ ),
    .B1(\heichips25_sap3/_1274_ ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][1] ),
    .A2(\heichips25_sap3/_1270_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][1] ));
 sg13g2_nand4_1 \heichips25_sap3/_3781_  (.B(\heichips25_sap3/_1289_ ),
    .C(\heichips25_sap3/_1290_ ),
    .A(\heichips25_sap3/_1288_ ),
    .Y(\heichips25_sap3/_1292_ ),
    .D(\heichips25_sap3/_1291_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_3782_  (.B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][1] ),
    .C1(\heichips25_sap3/_1292_ ),
    .B1(\heichips25_sap3/_1281_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][1] ),
    .Y(\heichips25_sap3/_1293_ ),
    .A2(\heichips25_sap3/_1272_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_3783_  (.B2(\heichips25_sap3/_1293_ ),
    .C1(\heichips25_sap3/net339 ),
    .B1(\heichips25_sap3/_1287_ ),
    .A1(\heichips25_sap3/_1385_ ),
    .Y(\heichips25_sap3/_1294_ ),
    .A2(\heichips25_sap3/net290 ));
 sg13g2_a21o_1 \heichips25_sap3/_3784_  (.A2(\heichips25_sap3/net339 ),
    .A1(\heichips25_sap3/net1141 ),
    .B1(\heichips25_sap3/_1294_ ),
    .X(\heichips25_sap3/_0174_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3785_  (.Y(\heichips25_sap3/_1295_ ),
    .B1(\heichips25_sap3/_1281_ ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][2] ),
    .A2(\heichips25_sap3/_1272_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][2] ));
 sg13g2_a22oi_1 \heichips25_sap3/_3786_  (.Y(\heichips25_sap3/_1296_ ),
    .B1(\heichips25_sap3/_1282_ ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][2] ),
    .A2(\heichips25_sap3/net292 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][2] ));
 sg13g2_a22oi_1 \heichips25_sap3/_3787_  (.Y(\heichips25_sap3/_1297_ ),
    .B1(\heichips25_sap3/_1279_ ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][2] ),
    .A2(\heichips25_sap3/_1278_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][2] ));
 sg13g2_a21oi_1 \heichips25_sap3/_3788_  (.A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][2] ),
    .A2(\heichips25_sap3/_1274_ ),
    .Y(\heichips25_sap3/_1298_ ),
    .B1(\heichips25_sap3/net290 ));
 sg13g2_a22oi_1 \heichips25_sap3/_3789_  (.Y(\heichips25_sap3/_1299_ ),
    .B1(\heichips25_sap3/net293 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][2] ),
    .A2(\heichips25_sap3/_1259_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][2] ));
 sg13g2_nand4_1 \heichips25_sap3/_3790_  (.B(\heichips25_sap3/_1296_ ),
    .C(\heichips25_sap3/_1298_ ),
    .A(\heichips25_sap3/_1295_ ),
    .Y(\heichips25_sap3/_1300_ ),
    .D(\heichips25_sap3/_1299_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_3791_  (.B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][2] ),
    .C1(\heichips25_sap3/_1300_ ),
    .B1(\heichips25_sap3/_1270_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][2] ),
    .Y(\heichips25_sap3/_1301_ ),
    .A2(\heichips25_sap3/_1265_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_3792_  (.B2(\heichips25_sap3/_1301_ ),
    .C1(\heichips25_sap3/net339 ),
    .B1(\heichips25_sap3/_1297_ ),
    .A1(\heichips25_sap3/_1375_ ),
    .Y(\heichips25_sap3/_1302_ ),
    .A2(\heichips25_sap3/net290 ));
 sg13g2_a21o_1 \heichips25_sap3/_3793_  (.A2(\heichips25_sap3/net339 ),
    .A1(\heichips25_sap3/net1120 ),
    .B1(\heichips25_sap3/_1302_ ),
    .X(\heichips25_sap3/_0175_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3794_  (.Y(\heichips25_sap3/_1303_ ),
    .B1(\heichips25_sap3/_1281_ ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][3] ),
    .A2(\heichips25_sap3/_1270_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][3] ));
 sg13g2_a22oi_1 \heichips25_sap3/_3795_  (.Y(\heichips25_sap3/_1304_ ),
    .B1(\heichips25_sap3/_1282_ ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][3] ),
    .A2(\heichips25_sap3/net292 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][3] ));
 sg13g2_a21oi_1 \heichips25_sap3/_3796_  (.A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][3] ),
    .A2(\heichips25_sap3/_1272_ ),
    .Y(\heichips25_sap3/_1305_ ),
    .B1(\heichips25_sap3/net290 ));
 sg13g2_a22oi_1 \heichips25_sap3/_3797_  (.Y(\heichips25_sap3/_1306_ ),
    .B1(\heichips25_sap3/_1279_ ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][3] ),
    .A2(\heichips25_sap3/net293 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][3] ));
 sg13g2_a22oi_1 \heichips25_sap3/_3798_  (.Y(\heichips25_sap3/_1307_ ),
    .B1(\heichips25_sap3/_1278_ ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][3] ),
    .A2(\heichips25_sap3/_1265_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][3] ));
 sg13g2_nand4_1 \heichips25_sap3/_3799_  (.B(\heichips25_sap3/_1305_ ),
    .C(\heichips25_sap3/_1306_ ),
    .A(\heichips25_sap3/_1304_ ),
    .Y(\heichips25_sap3/_1308_ ),
    .D(\heichips25_sap3/_1307_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_3800_  (.B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][3] ),
    .C1(\heichips25_sap3/_1308_ ),
    .B1(\heichips25_sap3/_1274_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][3] ),
    .Y(\heichips25_sap3/_1309_ ),
    .A2(\heichips25_sap3/_1259_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_3801_  (.B2(\heichips25_sap3/_1309_ ),
    .C1(\heichips25_sap3/net339 ),
    .B1(\heichips25_sap3/_1303_ ),
    .A1(\heichips25_sap3/_1368_ ),
    .Y(\heichips25_sap3/_1310_ ),
    .A2(\heichips25_sap3/net290 ));
 sg13g2_a21o_1 \heichips25_sap3/_3802_  (.A2(\heichips25_sap3/net340 ),
    .A1(\heichips25_sap3/net925 ),
    .B1(\heichips25_sap3/_1310_ ),
    .X(\heichips25_sap3/_0176_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3803_  (.Y(\heichips25_sap3/_1311_ ),
    .B1(\heichips25_sap3/_1282_ ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][4] ),
    .A2(\heichips25_sap3/_1270_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][4] ));
 sg13g2_a21oi_1 \heichips25_sap3/_3804_  (.A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][4] ),
    .A2(\heichips25_sap3/_1278_ ),
    .Y(\heichips25_sap3/_1312_ ),
    .B1(\heichips25_sap3/net291 ));
 sg13g2_a22oi_1 \heichips25_sap3/_3805_  (.Y(\heichips25_sap3/_1313_ ),
    .B1(\heichips25_sap3/_1281_ ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][4] ),
    .A2(\heichips25_sap3/_1259_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][4] ));
 sg13g2_a22oi_1 \heichips25_sap3/_3806_  (.Y(\heichips25_sap3/_1314_ ),
    .B1(\heichips25_sap3/_1279_ ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][4] ),
    .A2(\heichips25_sap3/net292 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][4] ));
 sg13g2_a22oi_1 \heichips25_sap3/_3807_  (.Y(\heichips25_sap3/_1315_ ),
    .B1(\heichips25_sap3/_1274_ ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][4] ),
    .A2(\heichips25_sap3/_1272_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][4] ));
 sg13g2_nand4_1 \heichips25_sap3/_3808_  (.B(\heichips25_sap3/_1313_ ),
    .C(\heichips25_sap3/_1314_ ),
    .A(\heichips25_sap3/_1312_ ),
    .Y(\heichips25_sap3/_1316_ ),
    .D(\heichips25_sap3/_1315_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_3809_  (.B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][4] ),
    .C1(\heichips25_sap3/_1316_ ),
    .B1(\heichips25_sap3/_1265_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][4] ),
    .Y(\heichips25_sap3/_1317_ ),
    .A2(\heichips25_sap3/net293 ));
 sg13g2_a221oi_1 \heichips25_sap3/_3810_  (.B2(\heichips25_sap3/_1317_ ),
    .C1(\heichips25_sap3/net340 ),
    .B1(\heichips25_sap3/_1311_ ),
    .A1(\heichips25_sap3/_1400_ ),
    .Y(\heichips25_sap3/_1318_ ),
    .A2(\heichips25_sap3/net291 ));
 sg13g2_a21o_1 \heichips25_sap3/_3811_  (.A2(\heichips25_sap3/net340 ),
    .A1(\heichips25_sap3/net891 ),
    .B1(\heichips25_sap3/_1318_ ),
    .X(\heichips25_sap3/_0177_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3812_  (.Y(\heichips25_sap3/_1319_ ),
    .B1(\heichips25_sap3/_1282_ ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][5] ),
    .A2(\heichips25_sap3/_1274_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][5] ));
 sg13g2_a22oi_1 \heichips25_sap3/_3813_  (.Y(\heichips25_sap3/_1320_ ),
    .B1(\heichips25_sap3/net292 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][5] ),
    .A2(\heichips25_sap3/_1265_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][5] ));
 sg13g2_a21oi_1 \heichips25_sap3/_3814_  (.A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][5] ),
    .A2(\heichips25_sap3/net293 ),
    .Y(\heichips25_sap3/_1321_ ),
    .B1(\heichips25_sap3/net291 ));
 sg13g2_a22oi_1 \heichips25_sap3/_3815_  (.Y(\heichips25_sap3/_1322_ ),
    .B1(\heichips25_sap3/_1281_ ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][5] ),
    .A2(\heichips25_sap3/_1279_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][5] ));
 sg13g2_a22oi_1 \heichips25_sap3/_3816_  (.Y(\heichips25_sap3/_1323_ ),
    .B1(\heichips25_sap3/_1278_ ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][5] ),
    .A2(\heichips25_sap3/_1272_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][5] ));
 sg13g2_nand4_1 \heichips25_sap3/_3817_  (.B(\heichips25_sap3/_1321_ ),
    .C(\heichips25_sap3/_1322_ ),
    .A(\heichips25_sap3/_1320_ ),
    .Y(\heichips25_sap3/_1324_ ),
    .D(\heichips25_sap3/_1323_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_3818_  (.B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][5] ),
    .C1(\heichips25_sap3/_1324_ ),
    .B1(\heichips25_sap3/_1270_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][5] ),
    .Y(\heichips25_sap3/_1325_ ),
    .A2(\heichips25_sap3/_1259_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_3819_  (.B2(\heichips25_sap3/_1325_ ),
    .C1(\heichips25_sap3/net340 ),
    .B1(\heichips25_sap3/_1319_ ),
    .A1(\heichips25_sap3/_1404_ ),
    .Y(\heichips25_sap3/_1326_ ),
    .A2(\heichips25_sap3/net291 ));
 sg13g2_a21o_1 \heichips25_sap3/_3820_  (.A2(\heichips25_sap3/net340 ),
    .A1(\heichips25_sap3/net1011 ),
    .B1(\heichips25_sap3/_1326_ ),
    .X(\heichips25_sap3/_0178_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3821_  (.A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][6] ),
    .A2(\heichips25_sap3/_1270_ ),
    .Y(\heichips25_sap3/_1327_ ),
    .B1(\heichips25_sap3/net291 ));
 sg13g2_a22oi_1 \heichips25_sap3/_3822_  (.Y(\heichips25_sap3/_1328_ ),
    .B1(\heichips25_sap3/net292 ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][6] ),
    .A2(\heichips25_sap3/_1259_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][6] ));
 sg13g2_a22oi_1 \heichips25_sap3/_3823_  (.Y(\heichips25_sap3/_1329_ ),
    .B1(\heichips25_sap3/_1279_ ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][6] ),
    .A2(\heichips25_sap3/_1274_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][6] ));
 sg13g2_a22oi_1 \heichips25_sap3/_3824_  (.Y(\heichips25_sap3/_1330_ ),
    .B1(\heichips25_sap3/_1281_ ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][6] ),
    .A2(\heichips25_sap3/_1272_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][6] ));
 sg13g2_a22oi_1 \heichips25_sap3/_3825_  (.Y(\heichips25_sap3/_1331_ ),
    .B1(\heichips25_sap3/_1265_ ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][6] ),
    .A2(\heichips25_sap3/net293 ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][6] ));
 sg13g2_nand4_1 \heichips25_sap3/_3826_  (.B(\heichips25_sap3/_1329_ ),
    .C(\heichips25_sap3/_1330_ ),
    .A(\heichips25_sap3/_1327_ ),
    .Y(\heichips25_sap3/_1332_ ),
    .D(\heichips25_sap3/_1331_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_3827_  (.B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][6] ),
    .C1(\heichips25_sap3/_1332_ ),
    .B1(\heichips25_sap3/_1282_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][6] ),
    .Y(\heichips25_sap3/_1333_ ),
    .A2(\heichips25_sap3/_1278_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_3828_  (.B2(\heichips25_sap3/_1333_ ),
    .C1(\heichips25_sap3/net340 ),
    .B1(\heichips25_sap3/_1328_ ),
    .A1(\heichips25_sap3/_1412_ ),
    .Y(\heichips25_sap3/_1334_ ),
    .A2(\heichips25_sap3/net291 ));
 sg13g2_a21o_1 \heichips25_sap3/_3829_  (.A2(\heichips25_sap3/net340 ),
    .A1(\heichips25_sap3/net953 ),
    .B1(\heichips25_sap3/_1334_ ),
    .X(\heichips25_sap3/_0179_ ));
 sg13g2_a22oi_1 \heichips25_sap3/_3830_  (.Y(\heichips25_sap3/_1335_ ),
    .B1(\heichips25_sap3/_1272_ ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][7] ),
    .A2(\heichips25_sap3/_1261_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][7] ));
 sg13g2_a22oi_1 \heichips25_sap3/_3831_  (.Y(\heichips25_sap3/_1336_ ),
    .B1(\heichips25_sap3/_1278_ ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][7] ),
    .A2(\heichips25_sap3/_1274_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][7] ));
 sg13g2_a22oi_1 \heichips25_sap3/_3832_  (.Y(\heichips25_sap3/_1337_ ),
    .B1(\heichips25_sap3/_1265_ ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][7] ),
    .A2(\heichips25_sap3/_1259_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][7] ));
 sg13g2_a21oi_1 \heichips25_sap3/_3833_  (.A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][7] ),
    .A2(\heichips25_sap3/_1279_ ),
    .Y(\heichips25_sap3/_1338_ ),
    .B1(\heichips25_sap3/net291 ));
 sg13g2_a22oi_1 \heichips25_sap3/_3834_  (.Y(\heichips25_sap3/_1339_ ),
    .B1(\heichips25_sap3/_1270_ ),
    .B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][7] ),
    .A2(\heichips25_sap3/_1266_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][7] ));
 sg13g2_nand4_1 \heichips25_sap3/_3835_  (.B(\heichips25_sap3/_1337_ ),
    .C(\heichips25_sap3/_1338_ ),
    .A(\heichips25_sap3/_1336_ ),
    .Y(\heichips25_sap3/_1340_ ),
    .D(\heichips25_sap3/_1339_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_3836_  (.B2(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][7] ),
    .C1(\heichips25_sap3/_1340_ ),
    .B1(\heichips25_sap3/_1282_ ),
    .A1(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][7] ),
    .Y(\heichips25_sap3/_1341_ ),
    .A2(\heichips25_sap3/_1281_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_3837_  (.B2(\heichips25_sap3/_1341_ ),
    .C1(\heichips25_sap3/_0008_ ),
    .B1(\heichips25_sap3/_1335_ ),
    .A1(\heichips25_sap3/_1420_ ),
    .Y(\heichips25_sap3/_1342_ ),
    .A2(\heichips25_sap3/net291 ));
 sg13g2_a21o_1 \heichips25_sap3/_3838_  (.A2(\heichips25_sap3/_0008_ ),
    .A1(\heichips25_sap3/net1031 ),
    .B1(\heichips25_sap3/_1342_ ),
    .X(\heichips25_sap3/_0180_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3839_  (.A(\heichips25_sap3/_1428_ ),
    .B(\heichips25_sap3/_0018_ ),
    .Y(\heichips25_sap3/_1343_ ));
 sg13g2_xnor2_1 \heichips25_sap3/_3840_  (.Y(\heichips25_sap3/_0181_ ),
    .A(\heichips25_sap3/net1197 ),
    .B(\heichips25_sap3/_0018_ ));
 sg13g2_xor2_1 \heichips25_sap3/_3841_  (.B(\heichips25_sap3/_1343_ ),
    .A(\heichips25_sap3/net1178 ),
    .X(\heichips25_sap3/_0182_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3842_  (.B1(\heichips25_sap3/net1224 ),
    .Y(\heichips25_sap3/_1344_ ),
    .A1(\heichips25_sap3/_0018_ ),
    .A2(\heichips25_sap3/_1260_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3843_  (.B1(\heichips25_sap3/_1344_ ),
    .Y(\heichips25_sap3/_0183_ ),
    .A1(\heichips25_sap3/_0018_ ),
    .A2(\heichips25_sap3/_1267_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3844_  (.B1(\heichips25_sap3/net1223 ),
    .Y(\heichips25_sap3/_1345_ ),
    .A1(\heichips25_sap3/_0018_ ),
    .A2(\heichips25_sap3/_1260_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3845_  (.B1(\heichips25_sap3/_1345_ ),
    .Y(\heichips25_sap3/_0184_ ),
    .A1(\heichips25_sap3/_0018_ ),
    .A2(\heichips25_sap3/_1262_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3846_  (.B1(\heichips25_sap3/_0288_ ),
    .Y(\heichips25_sap3/_1346_ ),
    .A1(\heichips25_sap3/net1225 ),
    .A2(\heichips25_sap3/_1366_ ));
 sg13g2_nor2_1 \heichips25_sap3/_3847_  (.A(\heichips25_sap3/net838 ),
    .B(\heichips25_sap3/_1346_ ),
    .Y(\heichips25_sap3/_1347_ ));
 sg13g2_mux4_1 \heichips25_sap3/_3848_  (.S0(\heichips25_sap3/net342 ),
    .A0(\heichips25_sap3/u_ser.shadow_reg[1] ),
    .A1(\heichips25_sap3/u_ser.shadow_reg[2] ),
    .A2(\heichips25_sap3/u_ser.shadow_reg[3] ),
    .A3(\heichips25_sap3/u_ser.shadow_reg[4] ),
    .S1(\heichips25_sap3/u_ser.bit_pos[1] ),
    .X(\heichips25_sap3/_1348_ ));
 sg13g2_nand3b_1 \heichips25_sap3/_3849_  (.B(\heichips25_sap3/u_ser.bit_pos[1] ),
    .C(\heichips25_sap3/u_ser.shadow_reg[7] ),
    .Y(\heichips25_sap3/_1349_ ),
    .A_N(\heichips25_sap3/net342 ));
 sg13g2_nand2b_1 \heichips25_sap3/_3850_  (.Y(\heichips25_sap3/_1350_ ),
    .B(\heichips25_sap3/net342 ),
    .A_N(\heichips25_sap3/u_ser.shadow_reg[6] ));
 sg13g2_o21ai_1 \heichips25_sap3/_3851_  (.B1(\heichips25_sap3/_1350_ ),
    .Y(\heichips25_sap3/_1351_ ),
    .A1(\heichips25_sap3/net342 ),
    .A2(\heichips25_sap3/u_ser.shadow_reg[5] ));
 sg13g2_o21ai_1 \heichips25_sap3/_3852_  (.B1(\heichips25_sap3/_1349_ ),
    .Y(\heichips25_sap3/_1352_ ),
    .A1(\heichips25_sap3/u_ser.bit_pos[1] ),
    .A2(\heichips25_sap3/_1351_ ));
 sg13g2_and3_1 \heichips25_sap3/_3853_  (.X(\heichips25_sap3/_1353_ ),
    .A(\heichips25_sap3/u_ser.state[1] ),
    .B(\heichips25_sap3/u_ser.bit_pos[2] ),
    .C(\heichips25_sap3/_1352_ ));
 sg13g2_a221oi_1 \heichips25_sap3/_3854_  (.B2(\heichips25_sap3/_1348_ ),
    .C1(\heichips25_sap3/_1353_ ),
    .B1(\heichips25_sap3/_0286_ ),
    .A1(\heichips25_sap3/_1359_ ),
    .Y(\heichips25_sap3/_1354_ ),
    .A2(\heichips25_sap3/u_ser.shadow_reg[0] ));
 sg13g2_a21oi_1 \heichips25_sap3/_3855_  (.A1(\heichips25_sap3/_1346_ ),
    .A2(\heichips25_sap3/_1354_ ),
    .Y(\heichips25_sap3/_0185_ ),
    .B1(\heichips25_sap3/_1347_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3856_  (.A1(\heichips25_sap3/_1430_ ),
    .A2(\heichips25_sap3/net341 ),
    .Y(\heichips25_sap3/_0186_ ),
    .B1(\heichips25_sap3/net830 ));
 sg13g2_nor2_1 \heichips25_sap3/_3857_  (.A(\heichips25_sap3/net1064 ),
    .B(\heichips25_sap3/net342 ),
    .Y(\heichips25_sap3/_1355_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3858_  (.A1(\heichips25_sap3/net342 ),
    .A2(\heichips25_sap3/_1346_ ),
    .Y(\heichips25_sap3/_0187_ ),
    .B1(\heichips25_sap3/_1355_ ));
 sg13g2_a21oi_1 \heichips25_sap3/_3859_  (.A1(\heichips25_sap3/net1071 ),
    .A2(\heichips25_sap3/_1346_ ),
    .Y(\heichips25_sap3/_1356_ ),
    .B1(\heichips25_sap3/u_ser.bit_pos[1] ));
 sg13g2_a21oi_1 \heichips25_sap3/_3860_  (.A1(\heichips25_sap3/net1065 ),
    .A2(\heichips25_sap3/_1346_ ),
    .Y(\heichips25_sap3/_0188_ ),
    .B1(\heichips25_sap3/net1072 ));
 sg13g2_o21ai_1 \heichips25_sap3/_3861_  (.B1(\heichips25_sap3/net1019 ),
    .Y(\heichips25_sap3/_1357_ ),
    .A1(\heichips25_sap3/net1064 ),
    .A2(\heichips25_sap3/_1366_ ));
 sg13g2_o21ai_1 \heichips25_sap3/_3862_  (.B1(\heichips25_sap3/_1357_ ),
    .Y(\heichips25_sap3/_0189_ ),
    .A1(\heichips25_sap3/_1359_ ),
    .A2(\heichips25_sap3/_1433_ ));
 sg13g2_mux2_1 \heichips25_sap3/_3863_  (.A0(\heichips25_sap3/sap_3_inst.out[0] ),
    .A1(\heichips25_sap3/net1145 ),
    .S(\heichips25_sap3/net341 ),
    .X(\heichips25_sap3/_0190_ ));
 sg13g2_mux2_1 \heichips25_sap3/_3864_  (.A0(\heichips25_sap3/sap_3_inst.out[1] ),
    .A1(\heichips25_sap3/net1121 ),
    .S(\heichips25_sap3/net341 ),
    .X(\heichips25_sap3/_0191_ ));
 sg13g2_mux2_1 \heichips25_sap3/_3865_  (.A0(\heichips25_sap3/sap_3_inst.out[2] ),
    .A1(\heichips25_sap3/net1149 ),
    .S(\heichips25_sap3/net341 ),
    .X(\heichips25_sap3/_0192_ ));
 sg13g2_mux2_1 \heichips25_sap3/_3866_  (.A0(\heichips25_sap3/sap_3_inst.out[3] ),
    .A1(\heichips25_sap3/net1119 ),
    .S(\heichips25_sap3/net341 ),
    .X(\heichips25_sap3/_0193_ ));
 sg13g2_mux2_1 \heichips25_sap3/_3867_  (.A0(\heichips25_sap3/sap_3_inst.out[4] ),
    .A1(\heichips25_sap3/net1143 ),
    .S(\heichips25_sap3/_0007_ ),
    .X(\heichips25_sap3/_0194_ ));
 sg13g2_mux2_1 \heichips25_sap3/_3868_  (.A0(\heichips25_sap3/sap_3_inst.out[5] ),
    .A1(\heichips25_sap3/net1124 ),
    .S(\heichips25_sap3/_0007_ ),
    .X(\heichips25_sap3/_0195_ ));
 sg13g2_mux2_1 \heichips25_sap3/_3869_  (.A0(\heichips25_sap3/sap_3_inst.out[6] ),
    .A1(\heichips25_sap3/net1105 ),
    .S(\heichips25_sap3/net341 ),
    .X(\heichips25_sap3/_0196_ ));
 sg13g2_mux2_1 \heichips25_sap3/_3870_  (.A0(\heichips25_sap3/sap_3_inst.out[7] ),
    .A1(\heichips25_sap3/net1112 ),
    .S(\heichips25_sap3/net341 ),
    .X(\heichips25_sap3/_0197_ ));
 sg13g2_inv_1 \heichips25_sap3/_3872__817  (.Y(net816),
    .A(\clknet_5_18__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_inv_1 \heichips25_sap3/_3873__818  (.Y(net817),
    .A(\clknet_5_16__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_inv_1 \heichips25_sap3/_3874__819  (.Y(net818),
    .A(\clknet_5_26__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_inv_1 \heichips25_sap3/_3875__820  (.Y(net819),
    .A(\clknet_5_27__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_inv_1 \heichips25_sap3/_3876__821  (.Y(net820),
    .A(\clknet_5_27__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_inv_1 \heichips25_sap3/_3877__822  (.Y(net821),
    .A(\clknet_5_27__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_inv_1 \heichips25_sap3/_3878__823  (.Y(net822),
    .A(\clknet_5_1__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_inv_1 \heichips25_sap3/_3879__824  (.Y(net823),
    .A(\clknet_5_1__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_inv_1 \heichips25_sap3/_3880__825  (.Y(net824),
    .A(\clknet_5_0__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_inv_1 \heichips25_sap3/_3881__826  (.Y(net825),
    .A(\clknet_5_0__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3882_  (.RESET_B(\heichips25_sap3/net450 ),
    .D(\heichips25_sap3/_0023_ ),
    .Q(\heichips25_sap3/sap_3_inst.out[0] ),
    .CLK(\clknet_5_17__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3883_  (.RESET_B(\heichips25_sap3/net450 ),
    .D(\heichips25_sap3/_0024_ ),
    .Q(\heichips25_sap3/sap_3_inst.out[1] ),
    .CLK(\clknet_5_17__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3884_  (.RESET_B(\heichips25_sap3/net450 ),
    .D(\heichips25_sap3/_0025_ ),
    .Q(\heichips25_sap3/sap_3_inst.out[2] ),
    .CLK(\clknet_5_17__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3885_  (.RESET_B(\heichips25_sap3/net451 ),
    .D(\heichips25_sap3/_0026_ ),
    .Q(\heichips25_sap3/sap_3_inst.out[3] ),
    .CLK(\clknet_5_20__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3886_  (.RESET_B(\heichips25_sap3/net453 ),
    .D(\heichips25_sap3/_0027_ ),
    .Q(\heichips25_sap3/sap_3_inst.out[4] ),
    .CLK(\clknet_5_21__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3887_  (.RESET_B(\heichips25_sap3/net451 ),
    .D(\heichips25_sap3/_0028_ ),
    .Q(\heichips25_sap3/sap_3_inst.out[5] ),
    .CLK(\clknet_5_20__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3888_  (.RESET_B(\heichips25_sap3/net451 ),
    .D(\heichips25_sap3/_0029_ ),
    .Q(\heichips25_sap3/sap_3_inst.out[6] ),
    .CLK(\clknet_5_20__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3889_  (.RESET_B(\heichips25_sap3/net451 ),
    .D(\heichips25_sap3/_0030_ ),
    .Q(\heichips25_sap3/sap_3_inst.out[7] ),
    .CLK(\clknet_5_20__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3890_  (.RESET_B(\heichips25_sap3/net447 ),
    .D(\heichips25_sap3/_0031_ ),
    .Q(\heichips25_sap3/sap_3_inst.alu_flags[2] ),
    .CLK(net814));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3891_  (.RESET_B(\heichips25_sap3/net447 ),
    .D(\heichips25_sap3/_0032_ ),
    .Q(\heichips25_sap3/sap_3_inst.alu_flags[3] ),
    .CLK(net815));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3892_  (.RESET_B(\heichips25_sap3/net435 ),
    .D(\heichips25_sap3/_0033_ ),
    .Q(\heichips25_sap3/sap_3_inst.alu_flags[0] ),
    .CLK(net816));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3893_  (.RESET_B(\heichips25_sap3/net435 ),
    .D(\heichips25_sap3/_0034_ ),
    .Q(\heichips25_sap3/sap_3_inst.alu_flags[1] ),
    .CLK(net817));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3894_  (.RESET_B(\heichips25_sap3/net448 ),
    .D(\heichips25_sap3/_0035_ ),
    .Q(\heichips25_sap3/sap_3_inst.alu_flags[4] ),
    .CLK(net818));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3895_  (.RESET_B(\heichips25_sap3/net448 ),
    .D(\heichips25_sap3/_0036_ ),
    .Q(\heichips25_sap3/sap_3_inst.alu_flags[5] ),
    .CLK(net819));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3896_  (.RESET_B(\heichips25_sap3/net448 ),
    .D(\heichips25_sap3/_0037_ ),
    .Q(\heichips25_sap3/sap_3_inst.alu_flags[6] ),
    .CLK(net820));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3897_  (.RESET_B(\heichips25_sap3/net449 ),
    .D(\heichips25_sap3/_0038_ ),
    .Q(\heichips25_sap3/sap_3_inst.alu_flags[7] ),
    .CLK(net821));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3898_  (.RESET_B(\heichips25_sap3/net450 ),
    .D(\heichips25_sap3/_0039_ ),
    .Q(\heichips25_sap3/sap_3_inst.alu_inst.carry ),
    .CLK(\clknet_5_16__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3899_  (.RESET_B(\heichips25_sap3/net447 ),
    .D(\heichips25_sap3/_0040_ ),
    .Q(\heichips25_sap3/sap_3_inst.alu_inst.acc[0] ),
    .CLK(\clknet_5_25__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3900_  (.RESET_B(\heichips25_sap3/net447 ),
    .D(\heichips25_sap3/_0041_ ),
    .Q(\heichips25_sap3/sap_3_inst.alu_inst.acc[1] ),
    .CLK(\clknet_5_26__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3901_  (.RESET_B(\heichips25_sap3/net448 ),
    .D(\heichips25_sap3/_0042_ ),
    .Q(\heichips25_sap3/sap_3_inst.alu_inst.acc[2] ),
    .CLK(\clknet_5_19__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3902_  (.RESET_B(\heichips25_sap3/net449 ),
    .D(\heichips25_sap3/_0043_ ),
    .Q(\heichips25_sap3/sap_3_inst.alu_inst.acc[3] ),
    .CLK(\clknet_5_22__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3903_  (.RESET_B(\heichips25_sap3/net455 ),
    .D(\heichips25_sap3/_0044_ ),
    .Q(\heichips25_sap3/sap_3_inst.alu_inst.acc[4] ),
    .CLK(\clknet_5_23__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3904_  (.RESET_B(\heichips25_sap3/net455 ),
    .D(\heichips25_sap3/_0045_ ),
    .Q(\heichips25_sap3/sap_3_inst.alu_inst.acc[5] ),
    .CLK(\clknet_5_23__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3905_  (.RESET_B(\heichips25_sap3/net455 ),
    .D(\heichips25_sap3/_0046_ ),
    .Q(\heichips25_sap3/sap_3_inst.alu_inst.acc[6] ),
    .CLK(\clknet_5_23__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3906_  (.RESET_B(\heichips25_sap3/net455 ),
    .D(\heichips25_sap3/_0047_ ),
    .Q(\heichips25_sap3/sap_3_inst.alu_inst.acc[7] ),
    .CLK(\clknet_5_22__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3907_  (.RESET_B(\heichips25_sap3/net447 ),
    .D(\heichips25_sap3/_0048_ ),
    .Q(\heichips25_sap3/sap_3_inst.alu_inst.act[0] ),
    .CLK(\clknet_5_18__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3908_  (.RESET_B(\heichips25_sap3/net447 ),
    .D(\heichips25_sap3/_0049_ ),
    .Q(\heichips25_sap3/sap_3_inst.alu_inst.act[1] ),
    .CLK(\clknet_5_27__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3909_  (.RESET_B(\heichips25_sap3/net448 ),
    .D(\heichips25_sap3/_0050_ ),
    .Q(\heichips25_sap3/sap_3_inst.alu_inst.act[2] ),
    .CLK(\clknet_5_19__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3910_  (.RESET_B(\heichips25_sap3/net448 ),
    .D(\heichips25_sap3/_0051_ ),
    .Q(\heichips25_sap3/sap_3_inst.alu_inst.act[3] ),
    .CLK(\clknet_5_19__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3911_  (.RESET_B(\heichips25_sap3/net455 ),
    .D(\heichips25_sap3/_0052_ ),
    .Q(\heichips25_sap3/sap_3_inst.alu_inst.act[4] ),
    .CLK(\clknet_5_21__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3912_  (.RESET_B(\heichips25_sap3/net454 ),
    .D(\heichips25_sap3/_0053_ ),
    .Q(\heichips25_sap3/sap_3_inst.alu_inst.act[5] ),
    .CLK(\clknet_5_21__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3913_  (.RESET_B(\heichips25_sap3/net454 ),
    .D(\heichips25_sap3/_0054_ ),
    .Q(\heichips25_sap3/sap_3_inst.alu_inst.act[6] ),
    .CLK(\clknet_5_21__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3914_  (.RESET_B(\heichips25_sap3/net455 ),
    .D(\heichips25_sap3/_0055_ ),
    .Q(\heichips25_sap3/sap_3_inst.alu_inst.act[7] ),
    .CLK(\clknet_5_23__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3915_  (.RESET_B(\heichips25_sap3/net450 ),
    .D(\heichips25_sap3/_0056_ ),
    .Q(\heichips25_sap3/sap_3_inst.alu_inst.tmp[0] ),
    .CLK(\clknet_5_17__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3916_  (.RESET_B(\heichips25_sap3/net435 ),
    .D(\heichips25_sap3/_0057_ ),
    .Q(\heichips25_sap3/sap_3_inst.alu_inst.tmp[1] ),
    .CLK(\clknet_5_18__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3917_  (.RESET_B(\heichips25_sap3/net447 ),
    .D(\heichips25_sap3/_0058_ ),
    .Q(\heichips25_sap3/sap_3_inst.alu_inst.tmp[2] ),
    .CLK(\clknet_5_19__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3918_  (.RESET_B(\heichips25_sap3/net449 ),
    .D(\heichips25_sap3/_0059_ ),
    .Q(\heichips25_sap3/sap_3_inst.alu_inst.tmp[3] ),
    .CLK(\clknet_5_22__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3919_  (.RESET_B(\heichips25_sap3/net448 ),
    .D(\heichips25_sap3/_0060_ ),
    .Q(\heichips25_sap3/sap_3_inst.alu_inst.tmp[4] ),
    .CLK(\clknet_5_22__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3920_  (.RESET_B(\heichips25_sap3/net448 ),
    .D(\heichips25_sap3/_0061_ ),
    .Q(\heichips25_sap3/sap_3_inst.alu_inst.tmp[5] ),
    .CLK(\clknet_5_22__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3921_  (.RESET_B(\heichips25_sap3/net450 ),
    .D(\heichips25_sap3/_0062_ ),
    .Q(\heichips25_sap3/sap_3_inst.alu_inst.tmp[6] ),
    .CLK(\clknet_5_20__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3922_  (.RESET_B(\heichips25_sap3/net450 ),
    .D(\heichips25_sap3/_0063_ ),
    .Q(\heichips25_sap3/sap_3_inst.alu_inst.tmp[7] ),
    .CLK(\clknet_5_17__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3923_  (.RESET_B(\heichips25_sap3/net435 ),
    .D(\heichips25_sap3/_0064_ ),
    .Q(\heichips25_sap3/sap_3_inst.controller_inst.opcode[0] ),
    .CLK(\clknet_5_16__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3924_  (.RESET_B(\heichips25_sap3/net435 ),
    .D(\heichips25_sap3/_0065_ ),
    .Q(\heichips25_sap3/sap_3_inst.controller_inst.opcode[1] ),
    .CLK(\clknet_5_24__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3925_  (.RESET_B(\heichips25_sap3/net435 ),
    .D(\heichips25_sap3/_0066_ ),
    .Q(\heichips25_sap3/sap_3_inst.controller_inst.opcode[2] ),
    .CLK(\clknet_5_5__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3926_  (.RESET_B(\heichips25_sap3/net436 ),
    .D(\heichips25_sap3/_0067_ ),
    .Q(\heichips25_sap3/sap_3_inst.controller_inst.opcode[3] ),
    .CLK(\clknet_5_18__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3927_  (.RESET_B(\heichips25_sap3/net436 ),
    .D(\heichips25_sap3/_0068_ ),
    .Q(\heichips25_sap3/sap_3_inst.controller_inst.opcode[4] ),
    .CLK(\clknet_5_18__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3928_  (.RESET_B(\heichips25_sap3/net436 ),
    .D(\heichips25_sap3/_0069_ ),
    .Q(\heichips25_sap3/sap_3_inst.controller_inst.opcode[5] ),
    .CLK(\clknet_5_5__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3929_  (.RESET_B(\heichips25_sap3/net435 ),
    .D(\heichips25_sap3/_0070_ ),
    .Q(\heichips25_sap3/sap_3_inst.controller_inst.opcode[6] ),
    .CLK(\clknet_5_16__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3930_  (.RESET_B(\heichips25_sap3/net435 ),
    .D(\heichips25_sap3/_0071_ ),
    .Q(\heichips25_sap3/sap_3_inst.controller_inst.opcode[7] ),
    .CLK(\clknet_5_16__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3931_  (.RESET_B(\heichips25_sap3/net438 ),
    .D(\heichips25_sap3/_0072_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[0][0] ),
    .CLK(\clknet_5_3__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3932_  (.RESET_B(\heichips25_sap3/net434 ),
    .D(\heichips25_sap3/_0073_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[0][1] ),
    .CLK(\clknet_5_4__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3933_  (.RESET_B(\heichips25_sap3/net433 ),
    .D(\heichips25_sap3/_0074_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[0][2] ),
    .CLK(\clknet_5_3__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3934_  (.RESET_B(\heichips25_sap3/net438 ),
    .D(\heichips25_sap3/_0075_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[0][3] ),
    .CLK(\clknet_5_2__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3935_  (.RESET_B(\heichips25_sap3/net438 ),
    .D(\heichips25_sap3/_0076_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[0][4] ),
    .CLK(\clknet_5_8__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3936_  (.RESET_B(\heichips25_sap3/net441 ),
    .D(\heichips25_sap3/_0077_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[0][5] ),
    .CLK(\clknet_5_10__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3937_  (.RESET_B(\heichips25_sap3/net441 ),
    .D(\heichips25_sap3/_0078_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[0][6] ),
    .CLK(\clknet_5_11__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3938_  (.RESET_B(\heichips25_sap3/net440 ),
    .D(\heichips25_sap3/_0079_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[0][7] ),
    .CLK(\clknet_5_9__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3939_  (.RESET_B(\heichips25_sap3/net456 ),
    .D(\heichips25_sap3/_0080_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][0] ),
    .CLK(\clknet_5_29__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3940_  (.RESET_B(\heichips25_sap3/net443 ),
    .D(\heichips25_sap3/_0081_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][1] ),
    .CLK(\clknet_5_5__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3941_  (.RESET_B(\heichips25_sap3/net456 ),
    .D(\heichips25_sap3/_0082_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][2] ),
    .CLK(\clknet_5_26__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3942_  (.RESET_B(\heichips25_sap3/net456 ),
    .D(\heichips25_sap3/_0083_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][3] ),
    .CLK(\clknet_5_29__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3943_  (.RESET_B(\heichips25_sap3/net444 ),
    .D(\heichips25_sap3/_0084_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][4] ),
    .CLK(\clknet_5_12__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3944_  (.RESET_B(\heichips25_sap3/net441 ),
    .D(\heichips25_sap3/_0085_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][5] ),
    .CLK(\clknet_5_14__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3945_  (.RESET_B(\heichips25_sap3/net444 ),
    .D(\heichips25_sap3/_0086_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][6] ),
    .CLK(\clknet_5_13__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3946_  (.RESET_B(\heichips25_sap3/net444 ),
    .D(\heichips25_sap3/_0087_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[1][7] ),
    .CLK(\clknet_5_14__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3947_  (.RESET_B(\heichips25_sap3/net439 ),
    .D(\heichips25_sap3/_0088_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][0] ),
    .CLK(\clknet_5_6__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3948_  (.RESET_B(\heichips25_sap3/net433 ),
    .D(\heichips25_sap3/_0089_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][1] ),
    .CLK(\clknet_5_1__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3949_  (.RESET_B(\heichips25_sap3/net433 ),
    .D(\heichips25_sap3/_0090_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][2] ),
    .CLK(\clknet_5_0__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3950_  (.RESET_B(\heichips25_sap3/net438 ),
    .D(\heichips25_sap3/_0091_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][3] ),
    .CLK(\clknet_5_2__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3951_  (.RESET_B(\heichips25_sap3/net439 ),
    .D(\heichips25_sap3/_0092_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][4] ),
    .CLK(\clknet_5_3__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3952_  (.RESET_B(\heichips25_sap3/net441 ),
    .D(\heichips25_sap3/_0093_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][5] ),
    .CLK(\clknet_5_11__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3953_  (.RESET_B(\heichips25_sap3/net440 ),
    .D(\heichips25_sap3/_0094_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][6] ),
    .CLK(\clknet_5_8__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3954_  (.RESET_B(\heichips25_sap3/net440 ),
    .D(\heichips25_sap3/_0095_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[2][7] ),
    .CLK(\clknet_5_10__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3955_  (.RESET_B(\heichips25_sap3/net456 ),
    .D(\heichips25_sap3/_0096_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][0] ),
    .CLK(\clknet_5_29__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3956_  (.RESET_B(\heichips25_sap3/net434 ),
    .D(\heichips25_sap3/_0097_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][1] ),
    .CLK(\clknet_5_4__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3957_  (.RESET_B(\heichips25_sap3/net436 ),
    .D(\heichips25_sap3/_0098_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][2] ),
    .CLK(\clknet_5_24__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3958_  (.RESET_B(\heichips25_sap3/net457 ),
    .D(\heichips25_sap3/_0099_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][3] ),
    .CLK(\clknet_5_28__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3959_  (.RESET_B(\heichips25_sap3/net459 ),
    .D(\heichips25_sap3/_0100_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][4] ),
    .CLK(\clknet_5_31__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3960_  (.RESET_B(\heichips25_sap3/net444 ),
    .D(\heichips25_sap3/_0101_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][5] ),
    .CLK(\clknet_5_15__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3961_  (.RESET_B(\heichips25_sap3/net459 ),
    .D(\heichips25_sap3/_0102_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][6] ),
    .CLK(\clknet_5_30__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3962_  (.RESET_B(\heichips25_sap3/net444 ),
    .D(\heichips25_sap3/_0103_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[3][7] ),
    .CLK(\clknet_5_14__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3963_  (.RESET_B(\heichips25_sap3/net443 ),
    .D(\heichips25_sap3/_0104_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][0] ),
    .CLK(\clknet_5_7__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3964_  (.RESET_B(\heichips25_sap3/net434 ),
    .D(\heichips25_sap3/_0105_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][1] ),
    .CLK(\clknet_5_1__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3965_  (.RESET_B(\heichips25_sap3/net433 ),
    .D(\heichips25_sap3/_0106_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][2] ),
    .CLK(\clknet_5_0__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3966_  (.RESET_B(\heichips25_sap3/net438 ),
    .D(\heichips25_sap3/_0107_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][3] ),
    .CLK(\clknet_5_2__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3967_  (.RESET_B(\heichips25_sap3/net443 ),
    .D(\heichips25_sap3/_0108_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][4] ),
    .CLK(\clknet_5_12__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3968_  (.RESET_B(\heichips25_sap3/net441 ),
    .D(\heichips25_sap3/_0109_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][5] ),
    .CLK(\clknet_5_10__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3969_  (.RESET_B(\heichips25_sap3/net440 ),
    .D(\heichips25_sap3/_0110_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][6] ),
    .CLK(\clknet_5_8__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3970_  (.RESET_B(\heichips25_sap3/net440 ),
    .D(\heichips25_sap3/_0111_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[4][7] ),
    .CLK(\clknet_5_9__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3971_  (.RESET_B(\heichips25_sap3/net456 ),
    .D(\heichips25_sap3/_0112_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][0] ),
    .CLK(\clknet_5_28__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3972_  (.RESET_B(\heichips25_sap3/net443 ),
    .D(\heichips25_sap3/_0113_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][1] ),
    .CLK(\clknet_5_5__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3973_  (.RESET_B(\heichips25_sap3/net447 ),
    .D(\heichips25_sap3/_0114_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][2] ),
    .CLK(\clknet_5_25__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3974_  (.RESET_B(\heichips25_sap3/net457 ),
    .D(\heichips25_sap3/_0115_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][3] ),
    .CLK(\clknet_5_28__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3975_  (.RESET_B(\heichips25_sap3/net459 ),
    .D(\heichips25_sap3/_0116_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][4] ),
    .CLK(\clknet_5_31__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3976_  (.RESET_B(\heichips25_sap3/net445 ),
    .D(\heichips25_sap3/_0117_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][5] ),
    .CLK(\clknet_5_30__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3977_  (.RESET_B(\heichips25_sap3/net459 ),
    .D(\heichips25_sap3/_0118_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][6] ),
    .CLK(\clknet_5_30__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3978_  (.RESET_B(\heichips25_sap3/net444 ),
    .D(\heichips25_sap3/_0119_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[5][7] ),
    .CLK(\clknet_5_13__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3979_  (.RESET_B(\heichips25_sap3/net443 ),
    .D(\heichips25_sap3/_0120_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][0] ),
    .CLK(\clknet_5_7__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3980_  (.RESET_B(\heichips25_sap3/net434 ),
    .D(\heichips25_sap3/_0121_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][1] ),
    .CLK(\clknet_5_4__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3981_  (.RESET_B(\heichips25_sap3/net434 ),
    .D(\heichips25_sap3/_0122_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][2] ),
    .CLK(\clknet_5_4__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3982_  (.RESET_B(\heichips25_sap3/net439 ),
    .D(\heichips25_sap3/_0123_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][3] ),
    .CLK(\clknet_5_6__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3983_  (.RESET_B(\heichips25_sap3/net439 ),
    .D(\heichips25_sap3/_0124_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][4] ),
    .CLK(\clknet_5_6__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3984_  (.RESET_B(\heichips25_sap3/net441 ),
    .D(\heichips25_sap3/_0125_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][5] ),
    .CLK(\clknet_5_11__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3985_  (.RESET_B(\heichips25_sap3/net441 ),
    .D(\heichips25_sap3/_0126_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][6] ),
    .CLK(\clknet_5_12__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3986_  (.RESET_B(\heichips25_sap3/net441 ),
    .D(\heichips25_sap3/_0127_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[6][7] ),
    .CLK(\clknet_5_11__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3987_  (.RESET_B(\heichips25_sap3/net457 ),
    .D(\heichips25_sap3/_0128_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][0] ),
    .CLK(\clknet_5_28__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3988_  (.RESET_B(\heichips25_sap3/net443 ),
    .D(\heichips25_sap3/_0129_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][1] ),
    .CLK(\clknet_5_5__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3989_  (.RESET_B(\heichips25_sap3/net456 ),
    .D(\heichips25_sap3/_0130_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][2] ),
    .CLK(\clknet_5_25__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3990_  (.RESET_B(\heichips25_sap3/net457 ),
    .D(\heichips25_sap3/_0131_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][3] ),
    .CLK(\clknet_5_28__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3991_  (.RESET_B(\heichips25_sap3/net459 ),
    .D(\heichips25_sap3/_0132_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][4] ),
    .CLK(\clknet_5_30__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3992_  (.RESET_B(\heichips25_sap3/net445 ),
    .D(\heichips25_sap3/_0133_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][5] ),
    .CLK(\clknet_5_15__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3993_  (.RESET_B(\heichips25_sap3/net459 ),
    .D(\heichips25_sap3/_0134_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][6] ),
    .CLK(\clknet_5_30__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3994_  (.RESET_B(\heichips25_sap3/net444 ),
    .D(\heichips25_sap3/_0135_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[7][7] ),
    .CLK(\clknet_5_14__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3995_  (.RESET_B(\heichips25_sap3/net439 ),
    .D(\heichips25_sap3/_0136_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][0] ),
    .CLK(\clknet_5_6__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3996_  (.RESET_B(\heichips25_sap3/net434 ),
    .D(\heichips25_sap3/_0137_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][1] ),
    .CLK(\clknet_5_1__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3997_  (.RESET_B(\heichips25_sap3/net438 ),
    .D(\heichips25_sap3/_0138_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][2] ),
    .CLK(\clknet_5_2__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3998_  (.RESET_B(\heichips25_sap3/net439 ),
    .D(\heichips25_sap3/_0139_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][3] ),
    .CLK(\clknet_5_3__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_3999_  (.RESET_B(\heichips25_sap3/net438 ),
    .D(\heichips25_sap3/_0140_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][4] ),
    .CLK(\clknet_5_8__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4000_  (.RESET_B(\heichips25_sap3/net440 ),
    .D(\heichips25_sap3/_0141_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][5] ),
    .CLK(\clknet_5_10__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4001_  (.RESET_B(\heichips25_sap3/net440 ),
    .D(\heichips25_sap3/_0142_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][6] ),
    .CLK(\clknet_5_9__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4002_  (.RESET_B(\heichips25_sap3/net442 ),
    .D(\heichips25_sap3/_0143_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[8][7] ),
    .CLK(\clknet_5_9__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4003_  (.RESET_B(\heichips25_sap3/net456 ),
    .D(\heichips25_sap3/_0144_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][0] ),
    .CLK(\clknet_5_25__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4004_  (.RESET_B(\heichips25_sap3/net436 ),
    .D(\heichips25_sap3/_0145_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][1] ),
    .CLK(\clknet_5_24__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4005_  (.RESET_B(\heichips25_sap3/net449 ),
    .D(\heichips25_sap3/_0146_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][2] ),
    .CLK(\clknet_5_24__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4006_  (.RESET_B(\heichips25_sap3/net443 ),
    .D(\heichips25_sap3/_0147_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][3] ),
    .CLK(\clknet_5_12__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4007_  (.RESET_B(\heichips25_sap3/net445 ),
    .D(\heichips25_sap3/_0148_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][4] ),
    .CLK(\clknet_5_13__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4008_  (.RESET_B(\heichips25_sap3/net445 ),
    .D(\heichips25_sap3/_0149_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][5] ),
    .CLK(\clknet_5_13__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4009_  (.RESET_B(\heichips25_sap3/net444 ),
    .D(\heichips25_sap3/_0150_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][6] ),
    .CLK(\clknet_5_12__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4010_  (.RESET_B(\heichips25_sap3/net445 ),
    .D(\heichips25_sap3/_0151_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[9][7] ),
    .CLK(\clknet_5_15__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4011_  (.RESET_B(\heichips25_sap3/net443 ),
    .D(\heichips25_sap3/_0152_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][0] ),
    .CLK(\clknet_5_7__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4012_  (.RESET_B(\heichips25_sap3/net434 ),
    .D(\heichips25_sap3/_0153_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][1] ),
    .CLK(\clknet_5_4__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4013_  (.RESET_B(\heichips25_sap3/net433 ),
    .D(\heichips25_sap3/_0154_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][2] ),
    .CLK(\clknet_5_0__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4014_  (.RESET_B(\heichips25_sap3/net438 ),
    .D(\heichips25_sap3/_0155_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][3] ),
    .CLK(\clknet_5_2__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4015_  (.RESET_B(\heichips25_sap3/net439 ),
    .D(\heichips25_sap3/_0156_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][4] ),
    .CLK(\clknet_5_6__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4016_  (.RESET_B(\heichips25_sap3/net442 ),
    .D(\heichips25_sap3/_0157_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][5] ),
    .CLK(\clknet_5_10__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4017_  (.RESET_B(\heichips25_sap3/net440 ),
    .D(\heichips25_sap3/_0158_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][6] ),
    .CLK(\clknet_5_8__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4018_  (.RESET_B(\heichips25_sap3/net442 ),
    .D(\heichips25_sap3/_0159_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[10][7] ),
    .CLK(\clknet_5_9__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4019_  (.RESET_B(\heichips25_sap3/net456 ),
    .D(\heichips25_sap3/_0160_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][0] ),
    .CLK(\clknet_5_26__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4020_  (.RESET_B(\heichips25_sap3/net446 ),
    .D(\heichips25_sap3/_0161_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][1] ),
    .CLK(\clknet_5_7__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4021_  (.RESET_B(\heichips25_sap3/net449 ),
    .D(\heichips25_sap3/_0162_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][2] ),
    .CLK(\clknet_5_26__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4022_  (.RESET_B(\heichips25_sap3/net457 ),
    .D(\heichips25_sap3/_0163_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][3] ),
    .CLK(\clknet_5_29__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4023_  (.RESET_B(\heichips25_sap3/net457 ),
    .D(\heichips25_sap3/_0164_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][4] ),
    .CLK(\clknet_5_31__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4024_  (.RESET_B(\heichips25_sap3/net442 ),
    .D(\heichips25_sap3/_0165_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][5] ),
    .CLK(\clknet_5_14__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4025_  (.RESET_B(\heichips25_sap3/net459 ),
    .D(\heichips25_sap3/_0166_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][6] ),
    .CLK(\clknet_5_31__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4026_  (.RESET_B(\heichips25_sap3/net445 ),
    .D(\heichips25_sap3/_0167_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.data[11][7] ),
    .CLK(\clknet_5_15__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4027_  (.RESET_B(\heichips25_sap3/net461 ),
    .D(\heichips25_sap3/net1059 ),
    .Q(\heichips25_sap3/regFile_serial ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4028_  (.RESET_B(\heichips25_sap3/net458 ),
    .D(\heichips25_sap3/net833 ),
    .Q(\heichips25_sap3/regFile_serial_start ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4029_  (.RESET_B(\heichips25_sap3/net461 ),
    .D(\heichips25_sap3/_0170_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos[0] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4030_  (.RESET_B(\heichips25_sap3/net461 ),
    .D(\heichips25_sap3/_0171_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos[1] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4031_  (.RESET_B(\heichips25_sap3/net461 ),
    .D(\heichips25_sap3/net837 ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos[2] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4032_  (.RESET_B(\heichips25_sap3/net458 ),
    .D(\heichips25_sap3/_0173_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[0] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4033_  (.RESET_B(\heichips25_sap3/net458 ),
    .D(\heichips25_sap3/_0174_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[1] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4034_  (.RESET_B(\heichips25_sap3/net458 ),
    .D(\heichips25_sap3/_0175_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[2] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4035_  (.RESET_B(\heichips25_sap3/net458 ),
    .D(\heichips25_sap3/net926 ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[3] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4036_  (.RESET_B(\heichips25_sap3/net461 ),
    .D(\heichips25_sap3/net892 ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[4] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4037_  (.RESET_B(\heichips25_sap3/net460 ),
    .D(\heichips25_sap3/net1012 ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[5] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4038_  (.RESET_B(\heichips25_sap3/net460 ),
    .D(\heichips25_sap3/net954 ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[6] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4039_  (.RESET_B(\heichips25_sap3/net461 ),
    .D(\heichips25_sap3/net1032 ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[7] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4040_  (.RESET_B(\heichips25_sap3/net462 ),
    .D(\heichips25_sap3/_0181_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.word_index[0] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4041_  (.RESET_B(\heichips25_sap3/net460 ),
    .D(\heichips25_sap3/net1179 ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.word_index[1] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4042_  (.RESET_B(\heichips25_sap3/net460 ),
    .D(\heichips25_sap3/_0183_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.word_index[2] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4043_  (.RESET_B(\heichips25_sap3/net460 ),
    .D(\heichips25_sap3/_0184_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.word_index[3] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4044_  (.RESET_B(\heichips25_sap3/net452 ),
    .D(\heichips25_sap3/net839 ),
    .Q(\heichips25_sap3/sap_3_outputReg_serial ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4045_  (.RESET_B(\heichips25_sap3/net453 ),
    .D(\heichips25_sap3/net831 ),
    .Q(\heichips25_sap3/sap_3_outputReg_start_sync ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4046_  (.RESET_B(\heichips25_sap3/net452 ),
    .D(\heichips25_sap3/_0187_ ),
    .Q(\heichips25_sap3/u_ser.bit_pos[0] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4047_  (.RESET_B(\heichips25_sap3/net452 ),
    .D(\heichips25_sap3/net1073 ),
    .Q(\heichips25_sap3/u_ser.bit_pos[1] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4048_  (.RESET_B(\heichips25_sap3/net452 ),
    .D(\heichips25_sap3/_0189_ ),
    .Q(\heichips25_sap3/u_ser.bit_pos[2] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4049_  (.RESET_B(\heichips25_sap3/net451 ),
    .D(\heichips25_sap3/_0190_ ),
    .Q(\heichips25_sap3/u_ser.shadow_reg[0] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4050_  (.RESET_B(\heichips25_sap3/net451 ),
    .D(\heichips25_sap3/_0191_ ),
    .Q(\heichips25_sap3/u_ser.shadow_reg[1] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4051_  (.RESET_B(\heichips25_sap3/net451 ),
    .D(\heichips25_sap3/_0192_ ),
    .Q(\heichips25_sap3/u_ser.shadow_reg[2] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4052_  (.RESET_B(\heichips25_sap3/net452 ),
    .D(\heichips25_sap3/_0193_ ),
    .Q(\heichips25_sap3/u_ser.shadow_reg[3] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4053_  (.RESET_B(\heichips25_sap3/net453 ),
    .D(\heichips25_sap3/net1144 ),
    .Q(\heichips25_sap3/u_ser.shadow_reg[4] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4054_  (.RESET_B(\heichips25_sap3/net452 ),
    .D(\heichips25_sap3/net1125 ),
    .Q(\heichips25_sap3/u_ser.shadow_reg[5] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4055_  (.RESET_B(\heichips25_sap3/net451 ),
    .D(\heichips25_sap3/_0196_ ),
    .Q(\heichips25_sap3/u_ser.shadow_reg[6] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4056_  (.RESET_B(\heichips25_sap3/net452 ),
    .D(\heichips25_sap3/_0197_ ),
    .Q(\heichips25_sap3/u_ser.shadow_reg[7] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4057_  (.RESET_B(\heichips25_sap3/net452 ),
    .D(\heichips25_sap3/net1020 ),
    .Q(\heichips25_sap3/_0007_ ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4058_  (.RESET_B(\heichips25_sap3/net453 ),
    .D(\heichips25_sap3/_0001_ ),
    .Q(\heichips25_sap3/u_ser.state[1] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4059_  (.RESET_B(\heichips25_sap3/net453 ),
    .D(\heichips25_sap3/u_ser.state[0] ),
    .Q(\heichips25_sap3/u_ser.state[2] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4060_  (.RESET_B(\heichips25_sap3/net462 ),
    .D(\heichips25_sap3/_0018_ ),
    .Q(\heichips25_sap3/_0008_ ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4061_  (.RESET_B(\heichips25_sap3/net459 ),
    .D(\heichips25_sap3/_0000_ ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.state[1] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4062_  (.RESET_B(\heichips25_sap3/net458 ),
    .D(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.state[0] ),
    .Q(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.state[2] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4063_  (.RESET_B(\heichips25_sap3/net433 ),
    .D(\heichips25_sap3/_0003_ ),
    .Q(\heichips25_sap3/sap_3_inst.controller_inst.stage[0] ),
    .CLK(net822));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4064_  (.RESET_B(\heichips25_sap3/net434 ),
    .D(\heichips25_sap3/_0004_ ),
    .Q(\heichips25_sap3/sap_3_inst.controller_inst.stage[1] ),
    .CLK(net823));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4065_  (.RESET_B(\heichips25_sap3/net433 ),
    .D(\heichips25_sap3/_0005_ ),
    .Q(\heichips25_sap3/sap_3_inst.controller_inst.stage[2] ),
    .CLK(net824));
 sg13g2_dfrbpq_1 \heichips25_sap3/_4066_  (.RESET_B(\heichips25_sap3/net433 ),
    .D(\heichips25_sap3/_0006_ ),
    .Q(\heichips25_sap3/sap_3_inst.controller_inst.stage[3] ),
    .CLK(net825));
 sg13g2_tielo _13__525 (.L_LO(net524));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_1 \heichips25_sap3/_4069_  (.A(\heichips25_sap3/mem_ram_we ),
    .X(\uo_out_sap3[0] ));
 sg13g2_buf_1 \heichips25_sap3/_4070_  (.A(\heichips25_sap3/mem_mar_we ),
    .X(\uo_out_sap3[1] ));
 sg13g2_buf_1 \heichips25_sap3/_4071_  (.A(\heichips25_sap3/sap_3_outputReg_serial ),
    .X(\uo_out_sap3[2] ));
 sg13g2_buf_1 \heichips25_sap3/_4072_  (.A(\heichips25_sap3/sap_3_outputReg_start_sync ),
    .X(\uo_out_sap3[3] ));
 sg13g2_buf_1 \heichips25_sap3/_4073_  (.A(\heichips25_sap3/regFile_serial ),
    .X(\uo_out_sap3[4] ));
 sg13g2_buf_1 \heichips25_sap3/_4074_  (.A(\heichips25_sap3/regFile_serial_start ),
    .X(\uo_out_sap3[5] ));
 sg13g2_inv_1 \heichips25_sap3/clk_div_param_inst/_1_  (.Y(\heichips25_sap3/clk_div_param_inst/_0_ ),
    .A(\heichips25_sap3/clk_div_param_inst/net834 ));
 sg13g2_dfrbpq_1 \heichips25_sap3/clk_div_param_inst/_2_  (.RESET_B(\heichips25_sap3/net450 ),
    .D(\heichips25_sap3/clk_div_param_inst/_0_ ),
    .Q(\heichips25_sap3/clk_div_param_inst/clk_out_reg ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_buf_16 \heichips25_sap3/clk_div_param_inst/clock_root  (.X(\heichips25_sap3/clk_div_out ),
    .A(\heichips25_sap3/clk_div_param_inst/clk_out_reg ));
 sg13g2_lgcp_1 \heichips25_sap3/sap_3_inst.clock.clock_gate_inst  (.GATE(\heichips25_sap3/_0002_ ),
    .CLK(\heichips25_sap3/clk_div_out ),
    .GCLK(\heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_1 input1 (.A(ena),
    .X(net1));
 sg13g2_buf_1 input2 (.A(rst_n),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[0]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[1]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[2]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[3]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[4]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[5]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(ui_in[6]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(ui_in[7]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[0]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[1]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[2]),
    .X(net13));
 sg13g2_buf_1 input14 (.A(uio_in[3]),
    .X(net14));
 sg13g2_buf_1 input15 (.A(uio_in[4]),
    .X(net15));
 sg13g2_buf_1 input16 (.A(uio_in[5]),
    .X(net16));
 sg13g2_buf_1 input17 (.A(uio_in[6]),
    .X(net17));
 sg13g2_buf_1 input18 (.A(uio_in[7]),
    .X(net18));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uio_oe[0]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uio_oe[1]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uio_oe[2]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uio_oe[3]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uio_oe[4]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uio_oe[5]));
 sg13g2_buf_1 output25 (.A(net25),
    .X(uio_oe[6]));
 sg13g2_buf_1 output26 (.A(net26),
    .X(uio_oe[7]));
 sg13g2_buf_1 output27 (.A(net27),
    .X(uio_out[0]));
 sg13g2_buf_1 output28 (.A(net28),
    .X(uio_out[1]));
 sg13g2_buf_1 output29 (.A(net29),
    .X(uio_out[2]));
 sg13g2_buf_1 output30 (.A(net30),
    .X(uio_out[3]));
 sg13g2_buf_1 output31 (.A(net31),
    .X(uio_out[4]));
 sg13g2_buf_1 output32 (.A(net32),
    .X(uio_out[5]));
 sg13g2_buf_1 output33 (.A(net33),
    .X(uio_out[6]));
 sg13g2_buf_1 output34 (.A(net34),
    .X(uio_out[7]));
 sg13g2_buf_1 output35 (.A(net35),
    .X(uo_out[0]));
 sg13g2_buf_1 output36 (.A(net36),
    .X(uo_out[1]));
 sg13g2_buf_1 output37 (.A(net37),
    .X(uo_out[2]));
 sg13g2_buf_1 output38 (.A(net38),
    .X(uo_out[3]));
 sg13g2_buf_1 output39 (.A(net39),
    .X(uo_out[4]));
 sg13g2_buf_1 output40 (.A(net40),
    .X(uo_out[5]));
 sg13g2_buf_1 output41 (.A(net41),
    .X(uo_out[6]));
 sg13g2_buf_1 output42 (.A(net42),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout43 (.A(\uio_out_sap3[6] ),
    .X(net43));
 sg13g2_buf_1 fanout44 (.A(\uio_out_sap3[2] ),
    .X(net44));
 sg13g2_buf_2 \heichips25_sap3/fanout45  (.A(\heichips25_sap3/_0242_ ),
    .X(\heichips25_sap3/net45 ));
 sg13g2_buf_2 fanout46 (.A(\uio_out_sap3[4] ),
    .X(net46));
 sg13g2_buf_4 fanout47 (.X(net47),
    .A(\uio_out_sap3[7] ));
 sg13g2_buf_1 \heichips25_sap3/fanout48  (.A(\heichips25_sap3/net49 ),
    .X(\heichips25_sap3/net48 ));
 sg13g2_buf_1 \heichips25_sap3/fanout49  (.A(\heichips25_sap3/_0871_ ),
    .X(\heichips25_sap3/net49 ));
 sg13g2_buf_1 \heichips25_sap3/fanout50  (.A(\heichips25_sap3/_0922_ ),
    .X(\heichips25_sap3/net50 ));
 sg13g2_buf_1 \heichips25_sap3/fanout51  (.A(\heichips25_sap3/_0898_ ),
    .X(\heichips25_sap3/net51 ));
 sg13g2_buf_1 \heichips25_sap3/fanout52  (.A(\heichips25_sap3/_0898_ ),
    .X(\heichips25_sap3/net52 ));
 sg13g2_buf_1 \heichips25_sap3/fanout53  (.A(\heichips25_sap3/_0786_ ),
    .X(\heichips25_sap3/net53 ));
 sg13g2_buf_1 \heichips25_sap3/fanout54  (.A(\heichips25_sap3/_0786_ ),
    .X(\heichips25_sap3/net54 ));
 sg13g2_buf_1 \heichips25_sap3/fanout55  (.A(\heichips25_sap3/_0748_ ),
    .X(\heichips25_sap3/net55 ));
 sg13g2_buf_1 \heichips25_sap3/fanout56  (.A(\heichips25_sap3/_1134_ ),
    .X(\heichips25_sap3/net56 ));
 sg13g2_buf_1 \heichips25_sap3/fanout57  (.A(\heichips25_sap3/net58 ),
    .X(\heichips25_sap3/net57 ));
 sg13g2_buf_1 \heichips25_sap3/fanout58  (.A(\heichips25_sap3/_1052_ ),
    .X(\heichips25_sap3/net58 ));
 sg13g2_buf_1 \heichips25_sap3/fanout59  (.A(\heichips25_sap3/_0830_ ),
    .X(\heichips25_sap3/net59 ));
 sg13g2_buf_1 \heichips25_sap3/fanout60  (.A(\heichips25_sap3/_0830_ ),
    .X(\heichips25_sap3/net60 ));
 sg13g2_buf_1 \heichips25_sap3/fanout61  (.A(\heichips25_sap3/net62 ),
    .X(\heichips25_sap3/net61 ));
 sg13g2_buf_1 \heichips25_sap3/fanout62  (.A(\heichips25_sap3/_0829_ ),
    .X(\heichips25_sap3/net62 ));
 sg13g2_buf_1 \heichips25_sap3/fanout63  (.A(\heichips25_sap3/_0810_ ),
    .X(\heichips25_sap3/net63 ));
 sg13g2_buf_1 \heichips25_sap3/fanout64  (.A(\heichips25_sap3/_0444_ ),
    .X(\heichips25_sap3/net64 ));
 sg13g2_buf_1 \heichips25_sap3/fanout65  (.A(\heichips25_sap3/_0444_ ),
    .X(\heichips25_sap3/net65 ));
 sg13g2_buf_1 \heichips25_sap3/fanout66  (.A(\heichips25_sap3/net67 ),
    .X(\heichips25_sap3/net66 ));
 sg13g2_buf_1 \heichips25_sap3/fanout67  (.A(\heichips25_sap3/_1593_ ),
    .X(\heichips25_sap3/net67 ));
 sg13g2_buf_1 \heichips25_sap3/fanout68  (.A(\heichips25_sap3/_0883_ ),
    .X(\heichips25_sap3/net68 ));
 sg13g2_buf_1 \heichips25_sap3/fanout69  (.A(\heichips25_sap3/net70 ),
    .X(\heichips25_sap3/net69 ));
 sg13g2_buf_1 \heichips25_sap3/fanout70  (.A(\heichips25_sap3/_0440_ ),
    .X(\heichips25_sap3/net70 ));
 sg13g2_buf_1 \heichips25_sap3/fanout71  (.A(\heichips25_sap3/_1746_ ),
    .X(\heichips25_sap3/net71 ));
 sg13g2_buf_1 \heichips25_sap3/fanout72  (.A(\heichips25_sap3/_1746_ ),
    .X(\heichips25_sap3/net72 ));
 sg13g2_buf_1 \heichips25_sap3/fanout73  (.A(\heichips25_sap3/net74 ),
    .X(\heichips25_sap3/net73 ));
 sg13g2_buf_2 \heichips25_sap3/fanout74  (.A(\heichips25_sap3/_1745_ ),
    .X(\heichips25_sap3/net74 ));
 sg13g2_buf_1 \heichips25_sap3/fanout75  (.A(\heichips25_sap3/net76 ),
    .X(\heichips25_sap3/net75 ));
 sg13g2_buf_1 \heichips25_sap3/fanout76  (.A(\heichips25_sap3/_1744_ ),
    .X(\heichips25_sap3/net76 ));
 sg13g2_buf_1 \heichips25_sap3/fanout77  (.A(\heichips25_sap3/net78 ),
    .X(\heichips25_sap3/net77 ));
 sg13g2_buf_1 \heichips25_sap3/fanout78  (.A(\heichips25_sap3/_1743_ ),
    .X(\heichips25_sap3/net78 ));
 sg13g2_buf_1 \heichips25_sap3/fanout79  (.A(\heichips25_sap3/_1741_ ),
    .X(\heichips25_sap3/net79 ));
 sg13g2_buf_1 \heichips25_sap3/fanout80  (.A(\heichips25_sap3/_1741_ ),
    .X(\heichips25_sap3/net80 ));
 sg13g2_buf_1 \heichips25_sap3/fanout81  (.A(\heichips25_sap3/net82 ),
    .X(\heichips25_sap3/net81 ));
 sg13g2_buf_1 \heichips25_sap3/fanout82  (.A(\heichips25_sap3/_1740_ ),
    .X(\heichips25_sap3/net82 ));
 sg13g2_buf_1 \heichips25_sap3/fanout83  (.A(\heichips25_sap3/_1739_ ),
    .X(\heichips25_sap3/net83 ));
 sg13g2_buf_1 \heichips25_sap3/fanout84  (.A(\heichips25_sap3/_1739_ ),
    .X(\heichips25_sap3/net84 ));
 sg13g2_buf_1 \heichips25_sap3/fanout85  (.A(\heichips25_sap3/net86 ),
    .X(\heichips25_sap3/net85 ));
 sg13g2_buf_1 \heichips25_sap3/fanout86  (.A(\heichips25_sap3/_1737_ ),
    .X(\heichips25_sap3/net86 ));
 sg13g2_buf_1 \heichips25_sap3/fanout87  (.A(\heichips25_sap3/net88 ),
    .X(\heichips25_sap3/net87 ));
 sg13g2_buf_1 \heichips25_sap3/fanout88  (.A(\heichips25_sap3/_1735_ ),
    .X(\heichips25_sap3/net88 ));
 sg13g2_buf_1 \heichips25_sap3/fanout89  (.A(\heichips25_sap3/net92 ),
    .X(\heichips25_sap3/net89 ));
 sg13g2_buf_1 \heichips25_sap3/fanout90  (.A(\heichips25_sap3/net92 ),
    .X(\heichips25_sap3/net90 ));
 sg13g2_buf_1 \heichips25_sap3/fanout91  (.A(\heichips25_sap3/net92 ),
    .X(\heichips25_sap3/net91 ));
 sg13g2_buf_1 \heichips25_sap3/fanout92  (.A(\heichips25_sap3/_1733_ ),
    .X(\heichips25_sap3/net92 ));
 sg13g2_buf_1 \heichips25_sap3/fanout93  (.A(\heichips25_sap3/_1187_ ),
    .X(\heichips25_sap3/net93 ));
 sg13g2_buf_1 \heichips25_sap3/fanout94  (.A(\heichips25_sap3/_1171_ ),
    .X(\heichips25_sap3/net94 ));
 sg13g2_buf_1 \heichips25_sap3/fanout95  (.A(\heichips25_sap3/_1144_ ),
    .X(\heichips25_sap3/net95 ));
 sg13g2_buf_1 \heichips25_sap3/fanout96  (.A(\heichips25_sap3/net97 ),
    .X(\heichips25_sap3/net96 ));
 sg13g2_buf_1 \heichips25_sap3/fanout97  (.A(\heichips25_sap3/net99 ),
    .X(\heichips25_sap3/net97 ));
 sg13g2_buf_1 \heichips25_sap3/fanout98  (.A(\heichips25_sap3/net99 ),
    .X(\heichips25_sap3/net98 ));
 sg13g2_buf_1 \heichips25_sap3/fanout99  (.A(\heichips25_sap3/_0862_ ),
    .X(\heichips25_sap3/net99 ));
 sg13g2_buf_1 \heichips25_sap3/fanout100  (.A(\heichips25_sap3/_0771_ ),
    .X(\heichips25_sap3/net100 ));
 sg13g2_buf_1 \heichips25_sap3/fanout101  (.A(\heichips25_sap3/_0771_ ),
    .X(\heichips25_sap3/net101 ));
 sg13g2_buf_1 \heichips25_sap3/fanout102  (.A(\heichips25_sap3/_0767_ ),
    .X(\heichips25_sap3/net102 ));
 sg13g2_buf_1 \heichips25_sap3/fanout103  (.A(\heichips25_sap3/_0767_ ),
    .X(\heichips25_sap3/net103 ));
 sg13g2_buf_1 \heichips25_sap3/fanout104  (.A(\heichips25_sap3/net105 ),
    .X(\heichips25_sap3/net104 ));
 sg13g2_buf_1 \heichips25_sap3/fanout105  (.A(\heichips25_sap3/_0763_ ),
    .X(\heichips25_sap3/net105 ));
 sg13g2_buf_1 \heichips25_sap3/fanout106  (.A(\heichips25_sap3/_0758_ ),
    .X(\heichips25_sap3/net106 ));
 sg13g2_buf_1 \heichips25_sap3/fanout107  (.A(\heichips25_sap3/_0758_ ),
    .X(\heichips25_sap3/net107 ));
 sg13g2_buf_1 \heichips25_sap3/fanout108  (.A(\heichips25_sap3/net110 ),
    .X(\heichips25_sap3/net108 ));
 sg13g2_buf_1 \heichips25_sap3/fanout109  (.A(\heichips25_sap3/net110 ),
    .X(\heichips25_sap3/net109 ));
 sg13g2_buf_1 \heichips25_sap3/fanout110  (.A(\heichips25_sap3/_0757_ ),
    .X(\heichips25_sap3/net110 ));
 sg13g2_buf_1 \heichips25_sap3/fanout111  (.A(\heichips25_sap3/net113 ),
    .X(\heichips25_sap3/net111 ));
 sg13g2_buf_1 \heichips25_sap3/fanout112  (.A(\heichips25_sap3/net113 ),
    .X(\heichips25_sap3/net112 ));
 sg13g2_buf_1 \heichips25_sap3/fanout113  (.A(\heichips25_sap3/_0755_ ),
    .X(\heichips25_sap3/net113 ));
 sg13g2_buf_1 \heichips25_sap3/fanout114  (.A(\heichips25_sap3/_0753_ ),
    .X(\heichips25_sap3/net114 ));
 sg13g2_buf_1 \heichips25_sap3/fanout115  (.A(\heichips25_sap3/_0753_ ),
    .X(\heichips25_sap3/net115 ));
 sg13g2_buf_1 \heichips25_sap3/fanout116  (.A(\heichips25_sap3/net118 ),
    .X(\heichips25_sap3/net116 ));
 sg13g2_buf_1 \heichips25_sap3/fanout117  (.A(\heichips25_sap3/net118 ),
    .X(\heichips25_sap3/net117 ));
 sg13g2_buf_1 \heichips25_sap3/fanout118  (.A(\heichips25_sap3/_0752_ ),
    .X(\heichips25_sap3/net118 ));
 sg13g2_buf_1 \heichips25_sap3/fanout119  (.A(\heichips25_sap3/_0750_ ),
    .X(\heichips25_sap3/net119 ));
 sg13g2_buf_1 \heichips25_sap3/fanout120  (.A(\heichips25_sap3/_0750_ ),
    .X(\heichips25_sap3/net120 ));
 sg13g2_buf_1 \heichips25_sap3/fanout121  (.A(\heichips25_sap3/net122 ),
    .X(\heichips25_sap3/net121 ));
 sg13g2_buf_1 \heichips25_sap3/fanout122  (.A(\heichips25_sap3/_0749_ ),
    .X(\heichips25_sap3/net122 ));
 sg13g2_buf_1 \heichips25_sap3/fanout123  (.A(\heichips25_sap3/_0720_ ),
    .X(\heichips25_sap3/net123 ));
 sg13g2_buf_1 \heichips25_sap3/fanout124  (.A(\heichips25_sap3/net126 ),
    .X(\heichips25_sap3/net124 ));
 sg13g2_buf_1 \heichips25_sap3/fanout125  (.A(\heichips25_sap3/net126 ),
    .X(\heichips25_sap3/net125 ));
 sg13g2_buf_1 \heichips25_sap3/fanout126  (.A(\heichips25_sap3/net130 ),
    .X(\heichips25_sap3/net126 ));
 sg13g2_buf_1 \heichips25_sap3/fanout127  (.A(\heichips25_sap3/net130 ),
    .X(\heichips25_sap3/net127 ));
 sg13g2_buf_1 \heichips25_sap3/fanout128  (.A(\heichips25_sap3/net130 ),
    .X(\heichips25_sap3/net128 ));
 sg13g2_buf_1 \heichips25_sap3/fanout129  (.A(\heichips25_sap3/net130 ),
    .X(\heichips25_sap3/net129 ));
 sg13g2_buf_1 \heichips25_sap3/fanout130  (.A(\heichips25_sap3/_0719_ ),
    .X(\heichips25_sap3/net130 ));
 sg13g2_buf_1 \heichips25_sap3/fanout131  (.A(\heichips25_sap3/_0881_ ),
    .X(\heichips25_sap3/net131 ));
 sg13g2_buf_1 \heichips25_sap3/fanout132  (.A(\heichips25_sap3/_0772_ ),
    .X(\heichips25_sap3/net132 ));
 sg13g2_buf_1 \heichips25_sap3/fanout133  (.A(\heichips25_sap3/_0772_ ),
    .X(\heichips25_sap3/net133 ));
 sg13g2_buf_1 \heichips25_sap3/fanout134  (.A(\heichips25_sap3/net137 ),
    .X(\heichips25_sap3/net134 ));
 sg13g2_buf_1 \heichips25_sap3/fanout135  (.A(\heichips25_sap3/net136 ),
    .X(\heichips25_sap3/net135 ));
 sg13g2_buf_1 \heichips25_sap3/fanout136  (.A(\heichips25_sap3/net137 ),
    .X(\heichips25_sap3/net136 ));
 sg13g2_buf_1 \heichips25_sap3/fanout137  (.A(\heichips25_sap3/_0770_ ),
    .X(\heichips25_sap3/net137 ));
 sg13g2_buf_1 \heichips25_sap3/fanout138  (.A(\heichips25_sap3/net139 ),
    .X(\heichips25_sap3/net138 ));
 sg13g2_buf_1 \heichips25_sap3/fanout139  (.A(\heichips25_sap3/_0768_ ),
    .X(\heichips25_sap3/net139 ));
 sg13g2_buf_1 \heichips25_sap3/fanout140  (.A(\heichips25_sap3/net141 ),
    .X(\heichips25_sap3/net140 ));
 sg13g2_buf_1 \heichips25_sap3/fanout141  (.A(\heichips25_sap3/net143 ),
    .X(\heichips25_sap3/net141 ));
 sg13g2_buf_1 \heichips25_sap3/fanout142  (.A(\heichips25_sap3/net143 ),
    .X(\heichips25_sap3/net142 ));
 sg13g2_buf_1 \heichips25_sap3/fanout143  (.A(\heichips25_sap3/_0766_ ),
    .X(\heichips25_sap3/net143 ));
 sg13g2_buf_1 \heichips25_sap3/fanout144  (.A(\heichips25_sap3/net145 ),
    .X(\heichips25_sap3/net144 ));
 sg13g2_buf_1 \heichips25_sap3/fanout145  (.A(\heichips25_sap3/_0760_ ),
    .X(\heichips25_sap3/net145 ));
 sg13g2_buf_1 \heichips25_sap3/fanout146  (.A(\heichips25_sap3/net149 ),
    .X(\heichips25_sap3/net146 ));
 sg13g2_buf_1 \heichips25_sap3/fanout147  (.A(\heichips25_sap3/net149 ),
    .X(\heichips25_sap3/net147 ));
 sg13g2_buf_1 \heichips25_sap3/fanout148  (.A(\heichips25_sap3/net149 ),
    .X(\heichips25_sap3/net148 ));
 sg13g2_buf_1 \heichips25_sap3/fanout149  (.A(\heichips25_sap3/_0754_ ),
    .X(\heichips25_sap3/net149 ));
 sg13g2_buf_1 \heichips25_sap3/fanout150  (.A(\heichips25_sap3/_0751_ ),
    .X(\heichips25_sap3/net150 ));
 sg13g2_buf_1 \heichips25_sap3/fanout151  (.A(\heichips25_sap3/_0751_ ),
    .X(\heichips25_sap3/net151 ));
 sg13g2_buf_1 \heichips25_sap3/fanout152  (.A(\heichips25_sap3/_0718_ ),
    .X(\heichips25_sap3/net152 ));
 sg13g2_buf_1 \heichips25_sap3/fanout153  (.A(\heichips25_sap3/_0606_ ),
    .X(\heichips25_sap3/net153 ));
 sg13g2_buf_1 \heichips25_sap3/fanout154  (.A(\heichips25_sap3/_0343_ ),
    .X(\heichips25_sap3/net154 ));
 sg13g2_buf_1 \heichips25_sap3/fanout155  (.A(\heichips25_sap3/net156 ),
    .X(\heichips25_sap3/net155 ));
 sg13g2_buf_1 \heichips25_sap3/fanout156  (.A(\heichips25_sap3/_1787_ ),
    .X(\heichips25_sap3/net156 ));
 sg13g2_buf_1 \heichips25_sap3/fanout157  (.A(\heichips25_sap3/net158 ),
    .X(\heichips25_sap3/net157 ));
 sg13g2_buf_1 \heichips25_sap3/fanout158  (.A(\heichips25_sap3/_0434_ ),
    .X(\heichips25_sap3/net158 ));
 sg13g2_buf_1 \heichips25_sap3/fanout159  (.A(\heichips25_sap3/_1895_ ),
    .X(\heichips25_sap3/net159 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout160  (.A(\heichips25_can_lehmann_fsm/net163 ),
    .X(\heichips25_can_lehmann_fsm/net160 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout161  (.A(\heichips25_can_lehmann_fsm/net163 ),
    .X(\heichips25_can_lehmann_fsm/net161 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout162  (.A(\heichips25_can_lehmann_fsm/net163 ),
    .X(\heichips25_can_lehmann_fsm/net162 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout163  (.A(\heichips25_can_lehmann_fsm/_0498_ ),
    .X(\heichips25_can_lehmann_fsm/net163 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout164  (.A(\heichips25_can_lehmann_fsm/net165 ),
    .X(\heichips25_can_lehmann_fsm/net164 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout165  (.A(\heichips25_can_lehmann_fsm/_0496_ ),
    .X(\heichips25_can_lehmann_fsm/net165 ));
 sg13g2_buf_1 \heichips25_sap3/fanout166  (.A(\heichips25_sap3/_0736_ ),
    .X(\heichips25_sap3/net166 ));
 sg13g2_buf_1 \heichips25_sap3/fanout167  (.A(\heichips25_sap3/_0605_ ),
    .X(\heichips25_sap3/net167 ));
 sg13g2_buf_1 \heichips25_sap3/fanout168  (.A(\heichips25_sap3/_1891_ ),
    .X(\heichips25_sap3/net168 ));
 sg13g2_buf_1 \heichips25_sap3/fanout169  (.A(\heichips25_sap3/_1891_ ),
    .X(\heichips25_sap3/net169 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout170  (.A(\heichips25_can_lehmann_fsm/net174 ),
    .X(\heichips25_can_lehmann_fsm/net170 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout171  (.A(\heichips25_can_lehmann_fsm/net173 ),
    .X(\heichips25_can_lehmann_fsm/net171 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout172  (.A(\heichips25_can_lehmann_fsm/net173 ),
    .X(\heichips25_can_lehmann_fsm/net172 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout173  (.A(\heichips25_can_lehmann_fsm/net174 ),
    .X(\heichips25_can_lehmann_fsm/net173 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout174  (.A(\heichips25_can_lehmann_fsm/_0557_ ),
    .X(\heichips25_can_lehmann_fsm/net174 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout175  (.A(\heichips25_can_lehmann_fsm/_0495_ ),
    .X(\heichips25_can_lehmann_fsm/net175 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout176  (.A(\heichips25_can_lehmann_fsm/_0495_ ),
    .X(\heichips25_can_lehmann_fsm/net176 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout177  (.A(\heichips25_can_lehmann_fsm/net180 ),
    .X(\heichips25_can_lehmann_fsm/net177 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout178  (.A(\heichips25_can_lehmann_fsm/net180 ),
    .X(\heichips25_can_lehmann_fsm/net178 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout179  (.A(\heichips25_can_lehmann_fsm/net180 ),
    .X(\heichips25_can_lehmann_fsm/net179 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout180  (.A(\heichips25_can_lehmann_fsm/_0313_ ),
    .X(\heichips25_can_lehmann_fsm/net180 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout181  (.A(\heichips25_can_lehmann_fsm/_0312_ ),
    .X(\heichips25_can_lehmann_fsm/net181 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout182  (.A(\heichips25_can_lehmann_fsm/net183 ),
    .X(\heichips25_can_lehmann_fsm/net182 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout183  (.A(\heichips25_can_lehmann_fsm/_0312_ ),
    .X(\heichips25_can_lehmann_fsm/net183 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout184  (.A(\heichips25_can_lehmann_fsm/net187 ),
    .X(\heichips25_can_lehmann_fsm/net184 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout185  (.A(\heichips25_can_lehmann_fsm/net187 ),
    .X(\heichips25_can_lehmann_fsm/net185 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout186  (.A(\heichips25_can_lehmann_fsm/net187 ),
    .X(\heichips25_can_lehmann_fsm/net186 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout187  (.A(\heichips25_can_lehmann_fsm/_0309_ ),
    .X(\heichips25_can_lehmann_fsm/net187 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout188  (.A(\heichips25_can_lehmann_fsm/net190 ),
    .X(\heichips25_can_lehmann_fsm/net188 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout189  (.A(\heichips25_can_lehmann_fsm/net190 ),
    .X(\heichips25_can_lehmann_fsm/net189 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout190  (.A(\heichips25_can_lehmann_fsm/_0307_ ),
    .X(\heichips25_can_lehmann_fsm/net190 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout191  (.A(\heichips25_can_lehmann_fsm/net192 ),
    .X(\heichips25_can_lehmann_fsm/net191 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout192  (.A(\heichips25_can_lehmann_fsm/net194 ),
    .X(\heichips25_can_lehmann_fsm/net192 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout193  (.A(\heichips25_can_lehmann_fsm/net194 ),
    .X(\heichips25_can_lehmann_fsm/net193 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout194  (.A(\heichips25_can_lehmann_fsm/_0306_ ),
    .X(\heichips25_can_lehmann_fsm/net194 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout195  (.A(\heichips25_can_lehmann_fsm/net196 ),
    .X(\heichips25_can_lehmann_fsm/net195 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout196  (.A(\heichips25_can_lehmann_fsm/_0306_ ),
    .X(\heichips25_can_lehmann_fsm/net196 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout197  (.A(\heichips25_can_lehmann_fsm/net200 ),
    .X(\heichips25_can_lehmann_fsm/net197 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout198  (.A(\heichips25_can_lehmann_fsm/net200 ),
    .X(\heichips25_can_lehmann_fsm/net198 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout199  (.A(\heichips25_can_lehmann_fsm/net200 ),
    .X(\heichips25_can_lehmann_fsm/net199 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout200  (.A(\heichips25_can_lehmann_fsm/_0305_ ),
    .X(\heichips25_can_lehmann_fsm/net200 ));
 sg13g2_buf_1 \heichips25_sap3/fanout201  (.A(\heichips25_sap3/_0624_ ),
    .X(\heichips25_sap3/net201 ));
 sg13g2_buf_1 \heichips25_sap3/fanout202  (.A(\heichips25_sap3/_0624_ ),
    .X(\heichips25_sap3/net202 ));
 sg13g2_buf_1 \heichips25_sap3/fanout203  (.A(\heichips25_sap3/net204 ),
    .X(\heichips25_sap3/net203 ));
 sg13g2_buf_1 \heichips25_sap3/fanout204  (.A(\heichips25_sap3/_0436_ ),
    .X(\heichips25_sap3/net204 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout205  (.A(\heichips25_can_lehmann_fsm/net210 ),
    .X(\heichips25_can_lehmann_fsm/net205 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout206  (.A(\heichips25_can_lehmann_fsm/net209 ),
    .X(\heichips25_can_lehmann_fsm/net206 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout207  (.A(\heichips25_can_lehmann_fsm/net208 ),
    .X(\heichips25_can_lehmann_fsm/net207 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout208  (.A(\heichips25_can_lehmann_fsm/net209 ),
    .X(\heichips25_can_lehmann_fsm/net208 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout209  (.A(\heichips25_can_lehmann_fsm/net210 ),
    .X(\heichips25_can_lehmann_fsm/net209 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout210  (.A(\heichips25_can_lehmann_fsm/_0476_ ),
    .X(\heichips25_can_lehmann_fsm/net210 ));
 sg13g2_buf_1 \heichips25_sap3/fanout211  (.A(\heichips25_sap3/net212 ),
    .X(\heichips25_sap3/net211 ));
 sg13g2_buf_1 \heichips25_sap3/fanout212  (.A(\heichips25_sap3/_1889_ ),
    .X(\heichips25_sap3/net212 ));
 sg13g2_buf_1 \heichips25_sap3/fanout213  (.A(\heichips25_sap3/net214 ),
    .X(\heichips25_sap3/net213 ));
 sg13g2_buf_1 \heichips25_sap3/fanout214  (.A(\heichips25_sap3/_0309_ ),
    .X(\heichips25_sap3/net214 ));
 sg13g2_buf_1 \heichips25_sap3/fanout215  (.A(\heichips25_sap3/_1801_ ),
    .X(\heichips25_sap3/net215 ));
 sg13g2_buf_1 \heichips25_sap3/fanout216  (.A(\heichips25_sap3/net218 ),
    .X(\heichips25_sap3/net216 ));
 sg13g2_buf_1 \heichips25_sap3/fanout217  (.A(\heichips25_sap3/net218 ),
    .X(\heichips25_sap3/net217 ));
 sg13g2_buf_1 \heichips25_sap3/fanout218  (.A(\heichips25_sap3/_1724_ ),
    .X(\heichips25_sap3/net218 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout219  (.A(\heichips25_can_lehmann_fsm/_1138_ ),
    .X(\heichips25_can_lehmann_fsm/net219 ));
 sg13g2_buf_1 \heichips25_sap3/fanout220  (.A(\heichips25_sap3/_1642_ ),
    .X(\heichips25_sap3/net220 ));
 sg13g2_buf_1 \heichips25_sap3/fanout221  (.A(\heichips25_sap3/_1642_ ),
    .X(\heichips25_sap3/net221 ));
 sg13g2_buf_1 \heichips25_sap3/fanout222  (.A(\heichips25_sap3/_1625_ ),
    .X(\heichips25_sap3/net222 ));
 sg13g2_buf_1 \heichips25_sap3/fanout223  (.A(\heichips25_sap3/_1622_ ),
    .X(\heichips25_sap3/net223 ));
 sg13g2_buf_1 \heichips25_sap3/fanout224  (.A(\heichips25_sap3/_1622_ ),
    .X(\heichips25_sap3/net224 ));
 sg13g2_buf_1 \heichips25_sap3/fanout225  (.A(\heichips25_sap3/_1598_ ),
    .X(\heichips25_sap3/net225 ));
 sg13g2_buf_1 \heichips25_sap3/fanout226  (.A(\heichips25_sap3/_1598_ ),
    .X(\heichips25_sap3/net226 ));
 sg13g2_buf_1 \heichips25_sap3/fanout227  (.A(\heichips25_sap3/net228 ),
    .X(\heichips25_sap3/net227 ));
 sg13g2_buf_1 \heichips25_sap3/fanout228  (.A(\heichips25_sap3/_1597_ ),
    .X(\heichips25_sap3/net228 ));
 sg13g2_buf_1 \heichips25_sap3/fanout229  (.A(\heichips25_sap3/_1497_ ),
    .X(\heichips25_sap3/net229 ));
 sg13g2_buf_1 \heichips25_sap3/fanout230  (.A(\heichips25_sap3/_1479_ ),
    .X(\heichips25_sap3/net230 ));
 sg13g2_buf_1 \heichips25_sap3/fanout231  (.A(\heichips25_sap3/net233 ),
    .X(\heichips25_sap3/net231 ));
 sg13g2_buf_1 \heichips25_sap3/fanout232  (.A(\heichips25_sap3/net233 ),
    .X(\heichips25_sap3/net232 ));
 sg13g2_buf_1 \heichips25_sap3/fanout233  (.A(\heichips25_sap3/_1466_ ),
    .X(\heichips25_sap3/net233 ));
 sg13g2_buf_1 \heichips25_sap3/fanout234  (.A(\heichips25_sap3/net235 ),
    .X(\heichips25_sap3/net234 ));
 sg13g2_buf_1 \heichips25_sap3/fanout235  (.A(\heichips25_sap3/_1462_ ),
    .X(\heichips25_sap3/net235 ));
 sg13g2_buf_1 \heichips25_sap3/fanout236  (.A(\heichips25_sap3/net240 ),
    .X(\heichips25_sap3/net236 ));
 sg13g2_buf_1 \heichips25_sap3/fanout237  (.A(\heichips25_sap3/net239 ),
    .X(\heichips25_sap3/net237 ));
 sg13g2_buf_1 \heichips25_sap3/fanout238  (.A(\heichips25_sap3/net239 ),
    .X(\heichips25_sap3/net238 ));
 sg13g2_buf_1 \heichips25_sap3/fanout239  (.A(\heichips25_sap3/net240 ),
    .X(\heichips25_sap3/net239 ));
 sg13g2_buf_1 \heichips25_sap3/fanout240  (.A(\heichips25_sap3/_1461_ ),
    .X(\heichips25_sap3/net240 ));
 sg13g2_buf_1 \heichips25_sap3/fanout241  (.A(\heichips25_sap3/_1452_ ),
    .X(\heichips25_sap3/net241 ));
 sg13g2_buf_1 \heichips25_sap3/fanout242  (.A(\heichips25_sap3/_1520_ ),
    .X(\heichips25_sap3/net242 ));
 sg13g2_buf_2 \heichips25_sap3/fanout243  (.A(\heichips25_sap3/_1512_ ),
    .X(\heichips25_sap3/net243 ));
 sg13g2_buf_1 \heichips25_sap3/fanout244  (.A(\heichips25_sap3/_1512_ ),
    .X(\heichips25_sap3/net244 ));
 sg13g2_buf_1 \heichips25_sap3/fanout245  (.A(\heichips25_sap3/_1509_ ),
    .X(\heichips25_sap3/net245 ));
 sg13g2_buf_1 \heichips25_sap3/fanout246  (.A(\heichips25_sap3/_1467_ ),
    .X(\heichips25_sap3/net246 ));
 sg13g2_buf_1 \heichips25_sap3/fanout247  (.A(\heichips25_sap3/_1457_ ),
    .X(\heichips25_sap3/net247 ));
 sg13g2_buf_1 \heichips25_sap3/fanout248  (.A(\heichips25_sap3/_1453_ ),
    .X(\heichips25_sap3/net248 ));
 sg13g2_buf_1 \heichips25_sap3/fanout249  (.A(\heichips25_sap3/_1451_ ),
    .X(\heichips25_sap3/net249 ));
 sg13g2_buf_1 \heichips25_sap3/fanout250  (.A(\heichips25_sap3/sap_3_inst.controller_inst.stage[3] ),
    .X(\heichips25_sap3/net250 ));
 sg13g2_buf_1 \heichips25_sap3/fanout251  (.A(\heichips25_sap3/sap_3_inst.controller_inst.stage[2] ),
    .X(\heichips25_sap3/net251 ));
 sg13g2_buf_1 \heichips25_sap3/fanout252  (.A(\heichips25_sap3/sap_3_inst.controller_inst.stage[1] ),
    .X(\heichips25_sap3/net252 ));
 sg13g2_buf_1 \heichips25_sap3/fanout253  (.A(\heichips25_sap3/sap_3_inst.controller_inst.stage[0] ),
    .X(\heichips25_sap3/net253 ));
 sg13g2_buf_1 \heichips25_sap3/fanout254  (.A(\heichips25_sap3/sap_3_inst.alu_flags[1] ),
    .X(\heichips25_sap3/net254 ));
 sg13g2_buf_1 \heichips25_sap3/fanout255  (.A(\heichips25_sap3/_1488_ ),
    .X(\heichips25_sap3/net255 ));
 sg13g2_buf_1 \heichips25_sap3/fanout256  (.A(\heichips25_sap3/_1442_ ),
    .X(\heichips25_sap3/net256 ));
 sg13g2_buf_1 \heichips25_sap3/fanout257  (.A(\heichips25_sap3/_1362_ ),
    .X(\heichips25_sap3/net257 ));
 sg13g2_buf_1 \heichips25_sap3/fanout258  (.A(\heichips25_sap3/sap_3_inst.controller_inst.opcode[7] ),
    .X(\heichips25_sap3/net258 ));
 sg13g2_buf_1 \heichips25_sap3/fanout259  (.A(\heichips25_sap3/sap_3_inst.controller_inst.opcode[7] ),
    .X(\heichips25_sap3/net259 ));
 sg13g2_buf_1 \heichips25_sap3/fanout260  (.A(\heichips25_sap3/sap_3_inst.controller_inst.opcode[6] ),
    .X(\heichips25_sap3/net260 ));
 sg13g2_buf_1 \heichips25_sap3/fanout261  (.A(\heichips25_sap3/sap_3_inst.controller_inst.opcode[5] ),
    .X(\heichips25_sap3/net261 ));
 sg13g2_buf_1 \heichips25_sap3/fanout262  (.A(\heichips25_sap3/net263 ),
    .X(\heichips25_sap3/net262 ));
 sg13g2_buf_1 \heichips25_sap3/fanout263  (.A(\heichips25_sap3/sap_3_inst.controller_inst.opcode[4] ),
    .X(\heichips25_sap3/net263 ));
 sg13g2_buf_1 \heichips25_sap3/fanout264  (.A(\heichips25_sap3/sap_3_inst.controller_inst.opcode[3] ),
    .X(\heichips25_sap3/net264 ));
 sg13g2_buf_1 \heichips25_sap3/fanout265  (.A(\heichips25_sap3/sap_3_inst.controller_inst.opcode[3] ),
    .X(\heichips25_sap3/net265 ));
 sg13g2_buf_1 \heichips25_sap3/fanout266  (.A(\heichips25_sap3/sap_3_inst.controller_inst.opcode[3] ),
    .X(\heichips25_sap3/net266 ));
 sg13g2_buf_1 \heichips25_sap3/fanout267  (.A(\heichips25_sap3/sap_3_inst.controller_inst.opcode[2] ),
    .X(\heichips25_sap3/net267 ));
 sg13g2_buf_1 \heichips25_sap3/fanout268  (.A(\heichips25_sap3/sap_3_inst.controller_inst.opcode[2] ),
    .X(\heichips25_sap3/net268 ));
 sg13g2_buf_1 \heichips25_sap3/fanout269  (.A(\heichips25_sap3/net270 ),
    .X(\heichips25_sap3/net269 ));
 sg13g2_buf_1 \heichips25_sap3/fanout270  (.A(\heichips25_sap3/net271 ),
    .X(\heichips25_sap3/net270 ));
 sg13g2_buf_1 \heichips25_sap3/fanout271  (.A(\heichips25_sap3/sap_3_inst.controller_inst.opcode[1] ),
    .X(\heichips25_sap3/net271 ));
 sg13g2_buf_1 \heichips25_sap3/fanout272  (.A(\heichips25_sap3/sap_3_inst.controller_inst.opcode[0] ),
    .X(\heichips25_sap3/net272 ));
 sg13g2_buf_1 \heichips25_sap3/fanout273  (.A(\heichips25_sap3/sap_3_inst.controller_inst.opcode[0] ),
    .X(\heichips25_sap3/net273 ));
 sg13g2_buf_1 \heichips25_sap3/fanout274  (.A(\heichips25_sap3/sap_3_inst.alu_inst.acc[7] ),
    .X(\heichips25_sap3/net274 ));
 sg13g2_buf_1 \heichips25_sap3/fanout275  (.A(\heichips25_sap3/sap_3_inst.alu_inst.acc[7] ),
    .X(\heichips25_sap3/net275 ));
 sg13g2_buf_1 \heichips25_sap3/fanout276  (.A(\heichips25_sap3/sap_3_inst.alu_inst.acc[6] ),
    .X(\heichips25_sap3/net276 ));
 sg13g2_buf_1 \heichips25_sap3/fanout277  (.A(\heichips25_sap3/sap_3_inst.alu_inst.acc[6] ),
    .X(\heichips25_sap3/net277 ));
 sg13g2_buf_1 \heichips25_sap3/fanout278  (.A(\heichips25_sap3/net279 ),
    .X(\heichips25_sap3/net278 ));
 sg13g2_buf_1 \heichips25_sap3/fanout279  (.A(\heichips25_sap3/sap_3_inst.alu_inst.acc[5] ),
    .X(\heichips25_sap3/net279 ));
 sg13g2_buf_1 \heichips25_sap3/fanout280  (.A(\heichips25_sap3/sap_3_inst.alu_inst.acc[4] ),
    .X(\heichips25_sap3/net280 ));
 sg13g2_buf_1 \heichips25_sap3/fanout281  (.A(\heichips25_sap3/sap_3_inst.alu_inst.acc[4] ),
    .X(\heichips25_sap3/net281 ));
 sg13g2_buf_1 \heichips25_sap3/fanout282  (.A(\heichips25_sap3/sap_3_inst.alu_inst.acc[3] ),
    .X(\heichips25_sap3/net282 ));
 sg13g2_buf_1 \heichips25_sap3/fanout283  (.A(\heichips25_sap3/sap_3_inst.alu_inst.acc[3] ),
    .X(\heichips25_sap3/net283 ));
 sg13g2_buf_1 \heichips25_sap3/fanout284  (.A(\heichips25_sap3/net285 ),
    .X(\heichips25_sap3/net284 ));
 sg13g2_buf_1 \heichips25_sap3/fanout285  (.A(\heichips25_sap3/sap_3_inst.alu_inst.acc[2] ),
    .X(\heichips25_sap3/net285 ));
 sg13g2_buf_1 \heichips25_sap3/fanout286  (.A(\heichips25_sap3/sap_3_inst.alu_inst.acc[1] ),
    .X(\heichips25_sap3/net286 ));
 sg13g2_buf_1 \heichips25_sap3/fanout287  (.A(\heichips25_sap3/sap_3_inst.alu_inst.acc[1] ),
    .X(\heichips25_sap3/net287 ));
 sg13g2_buf_1 \heichips25_sap3/fanout288  (.A(\heichips25_sap3/net289 ),
    .X(\heichips25_sap3/net288 ));
 sg13g2_buf_1 \heichips25_sap3/fanout289  (.A(\heichips25_sap3/sap_3_inst.alu_inst.acc[0] ),
    .X(\heichips25_sap3/net289 ));
 sg13g2_buf_1 \heichips25_sap3/fanout290  (.A(\heichips25_sap3/_1276_ ),
    .X(\heichips25_sap3/net290 ));
 sg13g2_buf_1 \heichips25_sap3/fanout291  (.A(\heichips25_sap3/_1276_ ),
    .X(\heichips25_sap3/net291 ));
 sg13g2_buf_1 \heichips25_sap3/fanout292  (.A(\heichips25_sap3/_1266_ ),
    .X(\heichips25_sap3/net292 ));
 sg13g2_buf_1 \heichips25_sap3/fanout293  (.A(\heichips25_sap3/_1261_ ),
    .X(\heichips25_sap3/net293 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout294  (.A(\heichips25_can_lehmann_fsm/_1004_ ),
    .X(\heichips25_can_lehmann_fsm/net294 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout295  (.A(\heichips25_can_lehmann_fsm/_1004_ ),
    .X(\heichips25_can_lehmann_fsm/net295 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout296  (.A(\heichips25_can_lehmann_fsm/net299 ),
    .X(\heichips25_can_lehmann_fsm/net296 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout297  (.A(\heichips25_can_lehmann_fsm/net299 ),
    .X(\heichips25_can_lehmann_fsm/net297 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout298  (.A(\heichips25_can_lehmann_fsm/net299 ),
    .X(\heichips25_can_lehmann_fsm/net298 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout299  (.A(\heichips25_can_lehmann_fsm/_1002_ ),
    .X(\heichips25_can_lehmann_fsm/net299 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout300  (.A(\heichips25_can_lehmann_fsm/net304 ),
    .X(\heichips25_can_lehmann_fsm/net300 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout301  (.A(\heichips25_can_lehmann_fsm/net304 ),
    .X(\heichips25_can_lehmann_fsm/net301 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout302  (.A(\heichips25_can_lehmann_fsm/net304 ),
    .X(\heichips25_can_lehmann_fsm/net302 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout303  (.A(\heichips25_can_lehmann_fsm/net304 ),
    .X(\heichips25_can_lehmann_fsm/net303 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout304  (.A(\heichips25_can_lehmann_fsm/_1000_ ),
    .X(\heichips25_can_lehmann_fsm/net304 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout305  (.A(\heichips25_can_lehmann_fsm/net309 ),
    .X(\heichips25_can_lehmann_fsm/net305 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout306  (.A(\heichips25_can_lehmann_fsm/net309 ),
    .X(\heichips25_can_lehmann_fsm/net306 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout307  (.A(\heichips25_can_lehmann_fsm/net309 ),
    .X(\heichips25_can_lehmann_fsm/net307 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout308  (.A(\heichips25_can_lehmann_fsm/net309 ),
    .X(\heichips25_can_lehmann_fsm/net308 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout309  (.A(\heichips25_can_lehmann_fsm/_0997_ ),
    .X(\heichips25_can_lehmann_fsm/net309 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout310  (.A(\heichips25_can_lehmann_fsm/net312 ),
    .X(\heichips25_can_lehmann_fsm/net310 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout311  (.A(\heichips25_can_lehmann_fsm/net312 ),
    .X(\heichips25_can_lehmann_fsm/net311 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout312  (.A(\heichips25_can_lehmann_fsm/_0994_ ),
    .X(\heichips25_can_lehmann_fsm/net312 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout313  (.A(\heichips25_can_lehmann_fsm/net316 ),
    .X(\heichips25_can_lehmann_fsm/net313 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout314  (.A(\heichips25_can_lehmann_fsm/net316 ),
    .X(\heichips25_can_lehmann_fsm/net314 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout315  (.A(\heichips25_can_lehmann_fsm/net316 ),
    .X(\heichips25_can_lehmann_fsm/net315 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout316  (.A(\heichips25_can_lehmann_fsm/_0993_ ),
    .X(\heichips25_can_lehmann_fsm/net316 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout317  (.A(\heichips25_can_lehmann_fsm/net320 ),
    .X(\heichips25_can_lehmann_fsm/net317 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout318  (.A(\heichips25_can_lehmann_fsm/net320 ),
    .X(\heichips25_can_lehmann_fsm/net318 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout319  (.A(\heichips25_can_lehmann_fsm/net320 ),
    .X(\heichips25_can_lehmann_fsm/net319 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout320  (.A(\heichips25_can_lehmann_fsm/_0990_ ),
    .X(\heichips25_can_lehmann_fsm/net320 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout321  (.A(\heichips25_can_lehmann_fsm/net324 ),
    .X(\heichips25_can_lehmann_fsm/net321 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout322  (.A(\heichips25_can_lehmann_fsm/net323 ),
    .X(\heichips25_can_lehmann_fsm/net322 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout323  (.A(\heichips25_can_lehmann_fsm/net324 ),
    .X(\heichips25_can_lehmann_fsm/net323 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout324  (.A(\heichips25_can_lehmann_fsm/net330 ),
    .X(\heichips25_can_lehmann_fsm/net324 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout325  (.A(\heichips25_can_lehmann_fsm/net326 ),
    .X(\heichips25_can_lehmann_fsm/net325 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout326  (.A(\heichips25_can_lehmann_fsm/net330 ),
    .X(\heichips25_can_lehmann_fsm/net326 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout327  (.A(\heichips25_can_lehmann_fsm/net329 ),
    .X(\heichips25_can_lehmann_fsm/net327 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout328  (.A(\heichips25_can_lehmann_fsm/net330 ),
    .X(\heichips25_can_lehmann_fsm/net328 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout329  (.A(\heichips25_can_lehmann_fsm/net330 ),
    .X(\heichips25_can_lehmann_fsm/net329 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout330  (.A(\heichips25_can_lehmann_fsm/_1175_ ),
    .X(\heichips25_can_lehmann_fsm/net330 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout331  (.A(\heichips25_can_lehmann_fsm/net334 ),
    .X(\heichips25_can_lehmann_fsm/net331 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout332  (.A(\heichips25_can_lehmann_fsm/net334 ),
    .X(\heichips25_can_lehmann_fsm/net332 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout333  (.A(\heichips25_can_lehmann_fsm/net334 ),
    .X(\heichips25_can_lehmann_fsm/net333 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout334  (.A(\heichips25_can_lehmann_fsm/_1003_ ),
    .X(\heichips25_can_lehmann_fsm/net334 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout335  (.A(\heichips25_can_lehmann_fsm/net336 ),
    .X(\heichips25_can_lehmann_fsm/net335 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout336  (.A(\heichips25_can_lehmann_fsm/_1001_ ),
    .X(\heichips25_can_lehmann_fsm/net336 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout337  (.A(\heichips25_can_lehmann_fsm/_0998_ ),
    .X(\heichips25_can_lehmann_fsm/net337 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout338  (.A(\heichips25_can_lehmann_fsm/_0983_ ),
    .X(\heichips25_can_lehmann_fsm/net338 ));
 sg13g2_buf_1 \heichips25_sap3/fanout339  (.A(\heichips25_sap3/net340 ),
    .X(\heichips25_sap3/net339 ));
 sg13g2_buf_1 \heichips25_sap3/fanout340  (.A(\heichips25_sap3/_0008_ ),
    .X(\heichips25_sap3/net340 ));
 sg13g2_buf_1 \heichips25_sap3/fanout341  (.A(\heichips25_sap3/net1276 ),
    .X(\heichips25_sap3/net341 ));
 sg13g2_buf_1 \heichips25_sap3/fanout342  (.A(\heichips25_sap3/net1071 ),
    .X(\heichips25_sap3/net342 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout343  (.A(\heichips25_can_lehmann_fsm/controller.extended_cond.opcode[0] ),
    .X(\heichips25_can_lehmann_fsm/net343 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout344  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[6] ),
    .X(\heichips25_can_lehmann_fsm/net344 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout345  (.A(\heichips25_can_lehmann_fsm/net1264 ),
    .X(\heichips25_can_lehmann_fsm/net345 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout346  (.A(\heichips25_can_lehmann_fsm/net1219 ),
    .X(\heichips25_can_lehmann_fsm/net346 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout347  (.A(\heichips25_can_lehmann_fsm/net1269 ),
    .X(\heichips25_can_lehmann_fsm/net347 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout348  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.addr[2] ),
    .X(\heichips25_can_lehmann_fsm/net348 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout349  (.A(\heichips25_can_lehmann_fsm/net350 ),
    .X(\heichips25_can_lehmann_fsm/net349 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout350  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.addr[2] ),
    .X(\heichips25_can_lehmann_fsm/net350 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout351  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.addr[1] ),
    .X(\heichips25_can_lehmann_fsm/net351 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout352  (.A(\heichips25_can_lehmann_fsm/net1273 ),
    .X(\heichips25_can_lehmann_fsm/net352 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout353  (.A(\heichips25_can_lehmann_fsm/net354 ),
    .X(\heichips25_can_lehmann_fsm/net353 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout354  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.addr[0] ),
    .X(\heichips25_can_lehmann_fsm/net354 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout355  (.A(\heichips25_can_lehmann_fsm/net356 ),
    .X(\heichips25_can_lehmann_fsm/net355 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout356  (.A(\heichips25_can_lehmann_fsm/net362 ),
    .X(\heichips25_can_lehmann_fsm/net356 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout357  (.A(\heichips25_can_lehmann_fsm/net358 ),
    .X(\heichips25_can_lehmann_fsm/net357 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout358  (.A(\heichips25_can_lehmann_fsm/net361 ),
    .X(\heichips25_can_lehmann_fsm/net358 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout359  (.A(\heichips25_can_lehmann_fsm/net360 ),
    .X(\heichips25_can_lehmann_fsm/net359 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout360  (.A(\heichips25_can_lehmann_fsm/net361 ),
    .X(\heichips25_can_lehmann_fsm/net360 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout361  (.A(\heichips25_can_lehmann_fsm/net362 ),
    .X(\heichips25_can_lehmann_fsm/net361 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout362  (.A(\heichips25_can_lehmann_fsm/net389 ),
    .X(\heichips25_can_lehmann_fsm/net362 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout363  (.A(\heichips25_can_lehmann_fsm/net364 ),
    .X(\heichips25_can_lehmann_fsm/net363 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout364  (.A(\heichips25_can_lehmann_fsm/net389 ),
    .X(\heichips25_can_lehmann_fsm/net364 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout365  (.A(\heichips25_can_lehmann_fsm/net367 ),
    .X(\heichips25_can_lehmann_fsm/net365 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout366  (.A(\heichips25_can_lehmann_fsm/net367 ),
    .X(\heichips25_can_lehmann_fsm/net366 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout367  (.A(\heichips25_can_lehmann_fsm/net389 ),
    .X(\heichips25_can_lehmann_fsm/net367 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout368  (.A(\heichips25_can_lehmann_fsm/net369 ),
    .X(\heichips25_can_lehmann_fsm/net368 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout369  (.A(\heichips25_can_lehmann_fsm/net371 ),
    .X(\heichips25_can_lehmann_fsm/net369 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout370  (.A(\heichips25_can_lehmann_fsm/net371 ),
    .X(\heichips25_can_lehmann_fsm/net370 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout371  (.A(\heichips25_can_lehmann_fsm/net373 ),
    .X(\heichips25_can_lehmann_fsm/net371 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout372  (.A(\heichips25_can_lehmann_fsm/net373 ),
    .X(\heichips25_can_lehmann_fsm/net372 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout373  (.A(\heichips25_can_lehmann_fsm/net389 ),
    .X(\heichips25_can_lehmann_fsm/net373 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout374  (.A(\heichips25_can_lehmann_fsm/net375 ),
    .X(\heichips25_can_lehmann_fsm/net374 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout375  (.A(\heichips25_can_lehmann_fsm/net379 ),
    .X(\heichips25_can_lehmann_fsm/net375 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout376  (.A(\heichips25_can_lehmann_fsm/net379 ),
    .X(\heichips25_can_lehmann_fsm/net376 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout377  (.A(\heichips25_can_lehmann_fsm/net379 ),
    .X(\heichips25_can_lehmann_fsm/net377 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout378  (.A(\heichips25_can_lehmann_fsm/net379 ),
    .X(\heichips25_can_lehmann_fsm/net378 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout379  (.A(\heichips25_can_lehmann_fsm/net389 ),
    .X(\heichips25_can_lehmann_fsm/net379 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout380  (.A(\heichips25_can_lehmann_fsm/net388 ),
    .X(\heichips25_can_lehmann_fsm/net380 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout381  (.A(\heichips25_can_lehmann_fsm/net388 ),
    .X(\heichips25_can_lehmann_fsm/net381 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout382  (.A(\heichips25_can_lehmann_fsm/net383 ),
    .X(\heichips25_can_lehmann_fsm/net382 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout383  (.A(\heichips25_can_lehmann_fsm/net388 ),
    .X(\heichips25_can_lehmann_fsm/net383 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout384  (.A(\heichips25_can_lehmann_fsm/net387 ),
    .X(\heichips25_can_lehmann_fsm/net384 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout385  (.A(\heichips25_can_lehmann_fsm/net387 ),
    .X(\heichips25_can_lehmann_fsm/net385 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout386  (.A(\heichips25_can_lehmann_fsm/net387 ),
    .X(\heichips25_can_lehmann_fsm/net386 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout387  (.A(\heichips25_can_lehmann_fsm/net388 ),
    .X(\heichips25_can_lehmann_fsm/net387 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout388  (.A(\heichips25_can_lehmann_fsm/net389 ),
    .X(\heichips25_can_lehmann_fsm/net388 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout389  (.A(\heichips25_can_lehmann_fsm/_0624_ ),
    .X(\heichips25_can_lehmann_fsm/net389 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout390  (.A(\heichips25_can_lehmann_fsm/net392 ),
    .X(\heichips25_can_lehmann_fsm/net390 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout391  (.A(\heichips25_can_lehmann_fsm/net392 ),
    .X(\heichips25_can_lehmann_fsm/net391 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout392  (.A(\heichips25_can_lehmann_fsm/net393 ),
    .X(\heichips25_can_lehmann_fsm/net392 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout393  (.A(\heichips25_can_lehmann_fsm/net408 ),
    .X(\heichips25_can_lehmann_fsm/net393 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout394  (.A(\heichips25_can_lehmann_fsm/net397 ),
    .X(\heichips25_can_lehmann_fsm/net394 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout395  (.A(\heichips25_can_lehmann_fsm/net397 ),
    .X(\heichips25_can_lehmann_fsm/net395 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout396  (.A(\heichips25_can_lehmann_fsm/net397 ),
    .X(\heichips25_can_lehmann_fsm/net396 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout397  (.A(\heichips25_can_lehmann_fsm/net400 ),
    .X(\heichips25_can_lehmann_fsm/net397 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout398  (.A(\heichips25_can_lehmann_fsm/net399 ),
    .X(\heichips25_can_lehmann_fsm/net398 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout399  (.A(\heichips25_can_lehmann_fsm/net400 ),
    .X(\heichips25_can_lehmann_fsm/net399 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout400  (.A(\heichips25_can_lehmann_fsm/net408 ),
    .X(\heichips25_can_lehmann_fsm/net400 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout401  (.A(\heichips25_can_lehmann_fsm/net402 ),
    .X(\heichips25_can_lehmann_fsm/net401 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout402  (.A(\heichips25_can_lehmann_fsm/net403 ),
    .X(\heichips25_can_lehmann_fsm/net402 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout403  (.A(\heichips25_can_lehmann_fsm/net408 ),
    .X(\heichips25_can_lehmann_fsm/net403 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout404  (.A(\heichips25_can_lehmann_fsm/net405 ),
    .X(\heichips25_can_lehmann_fsm/net404 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout405  (.A(\heichips25_can_lehmann_fsm/net407 ),
    .X(\heichips25_can_lehmann_fsm/net405 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout406  (.A(\heichips25_can_lehmann_fsm/net407 ),
    .X(\heichips25_can_lehmann_fsm/net406 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout407  (.A(\heichips25_can_lehmann_fsm/net408 ),
    .X(\heichips25_can_lehmann_fsm/net407 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout408  (.A(\heichips25_can_lehmann_fsm/net432 ),
    .X(\heichips25_can_lehmann_fsm/net408 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout409  (.A(\heichips25_can_lehmann_fsm/net411 ),
    .X(\heichips25_can_lehmann_fsm/net409 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout410  (.A(\heichips25_can_lehmann_fsm/net420 ),
    .X(\heichips25_can_lehmann_fsm/net410 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout411  (.A(\heichips25_can_lehmann_fsm/net420 ),
    .X(\heichips25_can_lehmann_fsm/net411 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout412  (.A(\heichips25_can_lehmann_fsm/net414 ),
    .X(\heichips25_can_lehmann_fsm/net412 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout413  (.A(\heichips25_can_lehmann_fsm/net414 ),
    .X(\heichips25_can_lehmann_fsm/net413 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout414  (.A(\heichips25_can_lehmann_fsm/net420 ),
    .X(\heichips25_can_lehmann_fsm/net414 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout415  (.A(\heichips25_can_lehmann_fsm/net416 ),
    .X(\heichips25_can_lehmann_fsm/net415 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout416  (.A(\heichips25_can_lehmann_fsm/net420 ),
    .X(\heichips25_can_lehmann_fsm/net416 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout417  (.A(\heichips25_can_lehmann_fsm/net419 ),
    .X(\heichips25_can_lehmann_fsm/net417 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout418  (.A(\heichips25_can_lehmann_fsm/net419 ),
    .X(\heichips25_can_lehmann_fsm/net418 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout419  (.A(\heichips25_can_lehmann_fsm/net420 ),
    .X(\heichips25_can_lehmann_fsm/net419 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout420  (.A(\heichips25_can_lehmann_fsm/net432 ),
    .X(\heichips25_can_lehmann_fsm/net420 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout421  (.A(\heichips25_can_lehmann_fsm/net422 ),
    .X(\heichips25_can_lehmann_fsm/net421 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout422  (.A(\heichips25_can_lehmann_fsm/net425 ),
    .X(\heichips25_can_lehmann_fsm/net422 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout423  (.A(\heichips25_can_lehmann_fsm/net425 ),
    .X(\heichips25_can_lehmann_fsm/net423 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout424  (.A(\heichips25_can_lehmann_fsm/net425 ),
    .X(\heichips25_can_lehmann_fsm/net424 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout425  (.A(\heichips25_can_lehmann_fsm/net432 ),
    .X(\heichips25_can_lehmann_fsm/net425 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout426  (.A(\heichips25_can_lehmann_fsm/net429 ),
    .X(\heichips25_can_lehmann_fsm/net426 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout427  (.A(\heichips25_can_lehmann_fsm/net429 ),
    .X(\heichips25_can_lehmann_fsm/net427 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout428  (.A(\heichips25_can_lehmann_fsm/net429 ),
    .X(\heichips25_can_lehmann_fsm/net428 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout429  (.A(\heichips25_can_lehmann_fsm/net431 ),
    .X(\heichips25_can_lehmann_fsm/net429 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout430  (.A(\heichips25_can_lehmann_fsm/net431 ),
    .X(\heichips25_can_lehmann_fsm/net430 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout431  (.A(\heichips25_can_lehmann_fsm/net432 ),
    .X(\heichips25_can_lehmann_fsm/net431 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout432  (.A(\heichips25_can_lehmann_fsm/_0623_ ),
    .X(\heichips25_can_lehmann_fsm/net432 ));
 sg13g2_buf_1 \heichips25_sap3/fanout433  (.A(\heichips25_sap3/net437 ),
    .X(\heichips25_sap3/net433 ));
 sg13g2_buf_1 \heichips25_sap3/fanout434  (.A(\heichips25_sap3/net437 ),
    .X(\heichips25_sap3/net434 ));
 sg13g2_buf_1 \heichips25_sap3/fanout435  (.A(\heichips25_sap3/net437 ),
    .X(\heichips25_sap3/net435 ));
 sg13g2_buf_1 \heichips25_sap3/fanout436  (.A(\heichips25_sap3/net437 ),
    .X(\heichips25_sap3/net436 ));
 sg13g2_buf_1 \heichips25_sap3/fanout437  (.A(_01_),
    .X(\heichips25_sap3/net437 ));
 sg13g2_buf_1 \heichips25_sap3/fanout438  (.A(\heichips25_sap3/net446 ),
    .X(\heichips25_sap3/net438 ));
 sg13g2_buf_1 \heichips25_sap3/fanout439  (.A(\heichips25_sap3/net446 ),
    .X(\heichips25_sap3/net439 ));
 sg13g2_buf_1 \heichips25_sap3/fanout440  (.A(\heichips25_sap3/net442 ),
    .X(\heichips25_sap3/net440 ));
 sg13g2_buf_1 \heichips25_sap3/fanout441  (.A(\heichips25_sap3/net442 ),
    .X(\heichips25_sap3/net441 ));
 sg13g2_buf_1 \heichips25_sap3/fanout442  (.A(\heichips25_sap3/net446 ),
    .X(\heichips25_sap3/net442 ));
 sg13g2_buf_1 \heichips25_sap3/fanout443  (.A(\heichips25_sap3/net446 ),
    .X(\heichips25_sap3/net443 ));
 sg13g2_buf_1 \heichips25_sap3/fanout444  (.A(\heichips25_sap3/net445 ),
    .X(\heichips25_sap3/net444 ));
 sg13g2_buf_1 \heichips25_sap3/fanout445  (.A(\heichips25_sap3/net446 ),
    .X(\heichips25_sap3/net445 ));
 sg13g2_buf_1 \heichips25_sap3/fanout446  (.A(_01_),
    .X(\heichips25_sap3/net446 ));
 sg13g2_buf_1 \heichips25_sap3/fanout447  (.A(\heichips25_sap3/net449 ),
    .X(\heichips25_sap3/net447 ));
 sg13g2_buf_1 \heichips25_sap3/fanout448  (.A(\heichips25_sap3/net449 ),
    .X(\heichips25_sap3/net448 ));
 sg13g2_buf_1 \heichips25_sap3/fanout449  (.A(\heichips25_sap3/net463 ),
    .X(\heichips25_sap3/net449 ));
 sg13g2_buf_1 \heichips25_sap3/fanout450  (.A(\heichips25_sap3/net463 ),
    .X(\heichips25_sap3/net450 ));
 sg13g2_buf_1 \heichips25_sap3/fanout451  (.A(\heichips25_sap3/net454 ),
    .X(\heichips25_sap3/net451 ));
 sg13g2_buf_1 \heichips25_sap3/fanout452  (.A(\heichips25_sap3/net453 ),
    .X(\heichips25_sap3/net452 ));
 sg13g2_buf_1 \heichips25_sap3/fanout453  (.A(\heichips25_sap3/net454 ),
    .X(\heichips25_sap3/net453 ));
 sg13g2_buf_1 \heichips25_sap3/fanout454  (.A(\heichips25_sap3/net455 ),
    .X(\heichips25_sap3/net454 ));
 sg13g2_buf_1 \heichips25_sap3/fanout455  (.A(\heichips25_sap3/net463 ),
    .X(\heichips25_sap3/net455 ));
 sg13g2_buf_1 \heichips25_sap3/fanout456  (.A(\heichips25_sap3/net458 ),
    .X(\heichips25_sap3/net456 ));
 sg13g2_buf_1 \heichips25_sap3/fanout457  (.A(\heichips25_sap3/net458 ),
    .X(\heichips25_sap3/net457 ));
 sg13g2_buf_1 \heichips25_sap3/fanout458  (.A(\heichips25_sap3/net462 ),
    .X(\heichips25_sap3/net458 ));
 sg13g2_buf_1 \heichips25_sap3/fanout459  (.A(\heichips25_sap3/net461 ),
    .X(\heichips25_sap3/net459 ));
 sg13g2_buf_1 \heichips25_sap3/fanout460  (.A(\heichips25_sap3/net461 ),
    .X(\heichips25_sap3/net460 ));
 sg13g2_buf_1 \heichips25_sap3/fanout461  (.A(\heichips25_sap3/net462 ),
    .X(\heichips25_sap3/net461 ));
 sg13g2_buf_1 \heichips25_sap3/fanout462  (.A(\heichips25_sap3/net463 ),
    .X(\heichips25_sap3/net462 ));
 sg13g2_buf_1 \heichips25_sap3/fanout463  (.A(_01_),
    .X(\heichips25_sap3/net463 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout464  (.A(\heichips25_can_lehmann_fsm/net466 ),
    .X(\heichips25_can_lehmann_fsm/net464 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout465  (.A(\heichips25_can_lehmann_fsm/net466 ),
    .X(\heichips25_can_lehmann_fsm/net465 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout466  (.A(\heichips25_can_lehmann_fsm/net470 ),
    .X(\heichips25_can_lehmann_fsm/net466 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout467  (.A(\heichips25_can_lehmann_fsm/net469 ),
    .X(\heichips25_can_lehmann_fsm/net467 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout468  (.A(\heichips25_can_lehmann_fsm/net469 ),
    .X(\heichips25_can_lehmann_fsm/net468 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout469  (.A(\heichips25_can_lehmann_fsm/net470 ),
    .X(\heichips25_can_lehmann_fsm/net469 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout470  (.A(\heichips25_can_lehmann_fsm/net503 ),
    .X(\heichips25_can_lehmann_fsm/net470 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout471  (.A(\heichips25_can_lehmann_fsm/net475 ),
    .X(\heichips25_can_lehmann_fsm/net471 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout472  (.A(\heichips25_can_lehmann_fsm/net474 ),
    .X(\heichips25_can_lehmann_fsm/net472 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout473  (.A(\heichips25_can_lehmann_fsm/net474 ),
    .X(\heichips25_can_lehmann_fsm/net473 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout474  (.A(\heichips25_can_lehmann_fsm/net475 ),
    .X(\heichips25_can_lehmann_fsm/net474 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout475  (.A(\heichips25_can_lehmann_fsm/net503 ),
    .X(\heichips25_can_lehmann_fsm/net475 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout476  (.A(\heichips25_can_lehmann_fsm/net479 ),
    .X(\heichips25_can_lehmann_fsm/net476 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout477  (.A(\heichips25_can_lehmann_fsm/net478 ),
    .X(\heichips25_can_lehmann_fsm/net477 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout478  (.A(\heichips25_can_lehmann_fsm/net479 ),
    .X(\heichips25_can_lehmann_fsm/net478 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout479  (.A(\heichips25_can_lehmann_fsm/net490 ),
    .X(\heichips25_can_lehmann_fsm/net479 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout480  (.A(\heichips25_can_lehmann_fsm/net481 ),
    .X(\heichips25_can_lehmann_fsm/net480 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout481  (.A(\heichips25_can_lehmann_fsm/net490 ),
    .X(\heichips25_can_lehmann_fsm/net481 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout482  (.A(\heichips25_can_lehmann_fsm/net484 ),
    .X(\heichips25_can_lehmann_fsm/net482 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout483  (.A(\heichips25_can_lehmann_fsm/net484 ),
    .X(\heichips25_can_lehmann_fsm/net483 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout484  (.A(\heichips25_can_lehmann_fsm/net490 ),
    .X(\heichips25_can_lehmann_fsm/net484 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout485  (.A(\heichips25_can_lehmann_fsm/net489 ),
    .X(\heichips25_can_lehmann_fsm/net485 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout486  (.A(\heichips25_can_lehmann_fsm/net489 ),
    .X(\heichips25_can_lehmann_fsm/net486 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout487  (.A(\heichips25_can_lehmann_fsm/net489 ),
    .X(\heichips25_can_lehmann_fsm/net487 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout488  (.A(\heichips25_can_lehmann_fsm/net489 ),
    .X(\heichips25_can_lehmann_fsm/net488 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout489  (.A(\heichips25_can_lehmann_fsm/net490 ),
    .X(\heichips25_can_lehmann_fsm/net489 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout490  (.A(\heichips25_can_lehmann_fsm/net503 ),
    .X(\heichips25_can_lehmann_fsm/net490 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout491  (.A(\heichips25_can_lehmann_fsm/net496 ),
    .X(\heichips25_can_lehmann_fsm/net491 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout492  (.A(\heichips25_can_lehmann_fsm/net493 ),
    .X(\heichips25_can_lehmann_fsm/net492 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout493  (.A(\heichips25_can_lehmann_fsm/net496 ),
    .X(\heichips25_can_lehmann_fsm/net493 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout494  (.A(\heichips25_can_lehmann_fsm/net496 ),
    .X(\heichips25_can_lehmann_fsm/net494 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout495  (.A(\heichips25_can_lehmann_fsm/net496 ),
    .X(\heichips25_can_lehmann_fsm/net495 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout496  (.A(\heichips25_can_lehmann_fsm/net503 ),
    .X(\heichips25_can_lehmann_fsm/net496 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout497  (.A(\heichips25_can_lehmann_fsm/net498 ),
    .X(\heichips25_can_lehmann_fsm/net497 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout498  (.A(\heichips25_can_lehmann_fsm/net502 ),
    .X(\heichips25_can_lehmann_fsm/net498 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout499  (.A(\heichips25_can_lehmann_fsm/net502 ),
    .X(\heichips25_can_lehmann_fsm/net499 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout500  (.A(\heichips25_can_lehmann_fsm/net502 ),
    .X(\heichips25_can_lehmann_fsm/net500 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout501  (.A(\heichips25_can_lehmann_fsm/net502 ),
    .X(\heichips25_can_lehmann_fsm/net501 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout502  (.A(\heichips25_can_lehmann_fsm/net503 ),
    .X(\heichips25_can_lehmann_fsm/net502 ));
 sg13g2_buf_1 \heichips25_can_lehmann_fsm/fanout503  (.A(_00_),
    .X(\heichips25_can_lehmann_fsm/net503 ));
 sg13g2_buf_1 fanout504 (.A(net506),
    .X(net504));
 sg13g2_buf_1 fanout505 (.A(net506),
    .X(net505));
 sg13g2_buf_1 fanout506 (.A(net1),
    .X(net506));
 sg13g2_buf_1 fanout507 (.A(net1),
    .X(net507));
 sg13g2_tielo _22__508 (.L_LO(net));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_16 clkbuf_0_clk (.X(clknet_0_clk),
    .A(clk));
 sg13g2_buf_16 clkbuf_2_0__f_clk (.X(clknet_2_0__leaf_clk),
    .A(clknet_0_clk));
 sg13g2_buf_16 clkbuf_2_1__f_clk (.X(clknet_2_1__leaf_clk),
    .A(clknet_0_clk));
 sg13g2_buf_16 clkbuf_2_2__f_clk (.X(clknet_2_2__leaf_clk),
    .A(clknet_0_clk));
 sg13g2_buf_16 clkbuf_2_3__f_clk (.X(clknet_2_3__leaf_clk),
    .A(clknet_0_clk));
 sg13g2_inv_4 clkload0 (.A(clknet_leaf_0_clk));
 sg13g2_inv_2 clkload1 (.A(clknet_leaf_1_clk));
 sg13g2_buf_8 clkload2 (.A(clknet_leaf_13_clk));
 sg13g2_inv_2 clkload3 (.A(clknet_leaf_21_clk));
 sg13g2_inv_2 clkload4 (.A(clknet_leaf_2_clk));
 sg13g2_inv_4 clkload5 (.A(clknet_leaf_3_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_leaf_4_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_leaf_5_clk));
 sg13g2_inv_2 clkload8 (.A(clknet_leaf_7_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_leaf_15_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_leaf_16_clk));
 sg13g2_buf_8 clkload11 (.A(clknet_leaf_17_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_leaf_20_clk));
 sg13g2_inv_2 clkload13 (.A(clknet_leaf_8_clk));
 sg13g2_buf_8 clkload14 (.A(clknet_leaf_9_clk));
 sg13g2_inv_2 clkload15 (.A(clknet_leaf_10_clk));
 sg13g2_inv_1 clkload16 (.A(clknet_leaf_11_clk));
 sg13g2_buf_8 clkload17 (.A(clknet_leaf_12_clk));
 sg13g2_buf_16 \clkbuf_0_heichips25_sap3/sap_3_inst.alu_inst.clk  (.X(\clknet_0_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .A(\heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_8 \clkbuf_4_0_0_heichips25_sap3/sap_3_inst.alu_inst.clk  (.A(\clknet_0_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .X(\clknet_4_0_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_8 \clkbuf_4_1_0_heichips25_sap3/sap_3_inst.alu_inst.clk  (.A(\clknet_0_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .X(\clknet_4_1_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_8 \clkbuf_4_2_0_heichips25_sap3/sap_3_inst.alu_inst.clk  (.A(\clknet_0_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .X(\clknet_4_2_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_8 \clkbuf_4_3_0_heichips25_sap3/sap_3_inst.alu_inst.clk  (.A(\clknet_0_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .X(\clknet_4_3_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_8 \clkbuf_4_4_0_heichips25_sap3/sap_3_inst.alu_inst.clk  (.A(\clknet_0_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .X(\clknet_4_4_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_8 \clkbuf_4_5_0_heichips25_sap3/sap_3_inst.alu_inst.clk  (.A(\clknet_0_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .X(\clknet_4_5_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_8 \clkbuf_4_6_0_heichips25_sap3/sap_3_inst.alu_inst.clk  (.A(\clknet_0_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .X(\clknet_4_6_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_8 \clkbuf_4_7_0_heichips25_sap3/sap_3_inst.alu_inst.clk  (.A(\clknet_0_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .X(\clknet_4_7_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_8 \clkbuf_4_8_0_heichips25_sap3/sap_3_inst.alu_inst.clk  (.A(\clknet_0_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .X(\clknet_4_8_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_8 \clkbuf_4_9_0_heichips25_sap3/sap_3_inst.alu_inst.clk  (.A(\clknet_0_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .X(\clknet_4_9_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_8 \clkbuf_4_10_0_heichips25_sap3/sap_3_inst.alu_inst.clk  (.A(\clknet_0_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .X(\clknet_4_10_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_8 \clkbuf_4_11_0_heichips25_sap3/sap_3_inst.alu_inst.clk  (.A(\clknet_0_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .X(\clknet_4_11_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_8 \clkbuf_4_12_0_heichips25_sap3/sap_3_inst.alu_inst.clk  (.A(\clknet_0_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .X(\clknet_4_12_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_8 \clkbuf_4_13_0_heichips25_sap3/sap_3_inst.alu_inst.clk  (.A(\clknet_0_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .X(\clknet_4_13_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_8 \clkbuf_4_14_0_heichips25_sap3/sap_3_inst.alu_inst.clk  (.A(\clknet_0_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .X(\clknet_4_14_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_8 \clkbuf_4_15_0_heichips25_sap3/sap_3_inst.alu_inst.clk  (.A(\clknet_0_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .X(\clknet_4_15_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_16 \clkbuf_5_0__f_heichips25_sap3/sap_3_inst.alu_inst.clk  (.X(\clknet_5_0__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .A(\clknet_4_0_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_16 \clkbuf_5_1__f_heichips25_sap3/sap_3_inst.alu_inst.clk  (.X(\clknet_5_1__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .A(\clknet_4_0_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_16 \clkbuf_5_2__f_heichips25_sap3/sap_3_inst.alu_inst.clk  (.X(\clknet_5_2__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .A(\clknet_4_1_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_16 \clkbuf_5_3__f_heichips25_sap3/sap_3_inst.alu_inst.clk  (.X(\clknet_5_3__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .A(\clknet_4_1_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_16 \clkbuf_5_4__f_heichips25_sap3/sap_3_inst.alu_inst.clk  (.X(\clknet_5_4__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .A(\clknet_4_2_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_16 \clkbuf_5_5__f_heichips25_sap3/sap_3_inst.alu_inst.clk  (.X(\clknet_5_5__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .A(\clknet_4_2_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_16 \clkbuf_5_6__f_heichips25_sap3/sap_3_inst.alu_inst.clk  (.X(\clknet_5_6__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .A(\clknet_4_3_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_16 \clkbuf_5_7__f_heichips25_sap3/sap_3_inst.alu_inst.clk  (.X(\clknet_5_7__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .A(\clknet_4_3_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_16 \clkbuf_5_8__f_heichips25_sap3/sap_3_inst.alu_inst.clk  (.X(\clknet_5_8__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .A(\clknet_4_4_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_16 \clkbuf_5_9__f_heichips25_sap3/sap_3_inst.alu_inst.clk  (.X(\clknet_5_9__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .A(\clknet_4_4_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_16 \clkbuf_5_10__f_heichips25_sap3/sap_3_inst.alu_inst.clk  (.X(\clknet_5_10__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .A(\clknet_4_5_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_16 \clkbuf_5_11__f_heichips25_sap3/sap_3_inst.alu_inst.clk  (.X(\clknet_5_11__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .A(\clknet_4_5_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_16 \clkbuf_5_12__f_heichips25_sap3/sap_3_inst.alu_inst.clk  (.X(\clknet_5_12__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .A(\clknet_4_6_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_16 \clkbuf_5_13__f_heichips25_sap3/sap_3_inst.alu_inst.clk  (.X(\clknet_5_13__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .A(\clknet_4_6_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_16 \clkbuf_5_14__f_heichips25_sap3/sap_3_inst.alu_inst.clk  (.X(\clknet_5_14__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .A(\clknet_4_7_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_16 \clkbuf_5_15__f_heichips25_sap3/sap_3_inst.alu_inst.clk  (.X(\clknet_5_15__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .A(\clknet_4_7_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_16 \clkbuf_5_16__f_heichips25_sap3/sap_3_inst.alu_inst.clk  (.X(\clknet_5_16__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .A(\clknet_4_8_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_16 \clkbuf_5_17__f_heichips25_sap3/sap_3_inst.alu_inst.clk  (.X(\clknet_5_17__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .A(\clknet_4_8_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_16 \clkbuf_5_18__f_heichips25_sap3/sap_3_inst.alu_inst.clk  (.X(\clknet_5_18__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .A(\clknet_4_9_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_16 \clkbuf_5_19__f_heichips25_sap3/sap_3_inst.alu_inst.clk  (.X(\clknet_5_19__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .A(\clknet_4_9_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_16 \clkbuf_5_20__f_heichips25_sap3/sap_3_inst.alu_inst.clk  (.X(\clknet_5_20__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .A(\clknet_4_10_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_16 \clkbuf_5_21__f_heichips25_sap3/sap_3_inst.alu_inst.clk  (.X(\clknet_5_21__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .A(\clknet_4_10_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_16 \clkbuf_5_22__f_heichips25_sap3/sap_3_inst.alu_inst.clk  (.X(\clknet_5_22__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .A(\clknet_4_11_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_16 \clkbuf_5_23__f_heichips25_sap3/sap_3_inst.alu_inst.clk  (.X(\clknet_5_23__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .A(\clknet_4_11_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_16 \clkbuf_5_24__f_heichips25_sap3/sap_3_inst.alu_inst.clk  (.X(\clknet_5_24__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .A(\clknet_4_12_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_16 \clkbuf_5_25__f_heichips25_sap3/sap_3_inst.alu_inst.clk  (.X(\clknet_5_25__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .A(\clknet_4_12_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_16 \clkbuf_5_26__f_heichips25_sap3/sap_3_inst.alu_inst.clk  (.X(\clknet_5_26__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .A(\clknet_4_13_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_16 \clkbuf_5_27__f_heichips25_sap3/sap_3_inst.alu_inst.clk  (.X(\clknet_5_27__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .A(\clknet_4_13_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_16 \clkbuf_5_28__f_heichips25_sap3/sap_3_inst.alu_inst.clk  (.X(\clknet_5_28__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .A(\clknet_4_14_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_16 \clkbuf_5_29__f_heichips25_sap3/sap_3_inst.alu_inst.clk  (.X(\clknet_5_29__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .A(\clknet_4_14_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_16 \clkbuf_5_30__f_heichips25_sap3/sap_3_inst.alu_inst.clk  (.X(\clknet_5_30__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .A(\clknet_4_15_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_16 \clkbuf_5_31__f_heichips25_sap3/sap_3_inst.alu_inst.clk  (.X(\clknet_5_31__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ),
    .A(\clknet_4_15_0_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_inv_1 clkload18 (.A(\clknet_5_3__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_inv_1 clkload19 (.A(\clknet_5_7__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_inv_1 clkload20 (.A(\clknet_5_11__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_inv_1 clkload21 (.A(\clknet_5_13__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_inv_1 clkload22 (.A(\clknet_5_15__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_inv_1 clkload23 (.A(\clknet_5_16__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_inv_1 clkload24 (.A(\clknet_5_19__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_inv_1 clkload25 (.A(\clknet_5_21__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_inv_1 clkload26 (.A(\clknet_5_23__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_inv_1 clkload27 (.A(\clknet_5_27__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_inv_1 clkload28 (.A(\clknet_5_29__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_inv_1 clkload29 (.A(\clknet_5_31__leaf_heichips25_sap3/sap_3_inst.alu_inst.clk ));
 sg13g2_buf_1 \heichips25_sap3/rebuffer827  (.A(\uio_out_sap3[6] ),
    .X(\heichips25_sap3/net826 ));
 sg13g2_buf_1 \heichips25_sap3/rebuffer828  (.A(\heichips25_sap3/_1736_ ),
    .X(\heichips25_sap3/net827 ));
 sg13g2_buf_1 \heichips25_sap3/rebuffer829  (.A(net829),
    .X(\heichips25_sap3/net828 ));
 sg13g2_buf_2 rebuffer830 (.A(\uio_oe_sap3[5] ),
    .X(net829));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold831  (.A(\heichips25_sap3/u_ser.state[2] ),
    .X(\heichips25_sap3/net830 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold832  (.A(\heichips25_sap3/_0186_ ),
    .X(\heichips25_sap3/net831 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold833  (.A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.state[2] ),
    .X(\heichips25_sap3/net832 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold834  (.A(\heichips25_sap3/_0169_ ),
    .X(\heichips25_sap3/net833 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/clk_div_param_inst/hold835  (.A(\heichips25_sap3/clk_div_param_inst/clk_out_reg ),
    .X(\heichips25_sap3/clk_div_param_inst/net834 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold836  (.A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos[2] ),
    .X(\heichips25_sap3/net835 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold837  (.A(\heichips25_sap3/_1256_ ),
    .X(\heichips25_sap3/net836 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold838  (.A(\heichips25_sap3/_0172_ ),
    .X(\heichips25_sap3/net837 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold839  (.A(\heichips25_sap3/sap_3_outputReg_serial ),
    .X(\heichips25_sap3/net838 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold840  (.A(\heichips25_sap3/_0185_ ),
    .X(\heichips25_sap3/net839 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold841  (.A(\heichips25_can_lehmann_fsm/controller.const_data[17] ),
    .X(\heichips25_can_lehmann_fsm/net840 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold842  (.A(\heichips25_can_lehmann_fsm/_0077_ ),
    .X(\heichips25_can_lehmann_fsm/net841 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold843  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[4] ),
    .X(\heichips25_can_lehmann_fsm/net842 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold844  (.A(\heichips25_can_lehmann_fsm/_0264_ ),
    .X(\heichips25_can_lehmann_fsm/net843 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold845  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[165] ),
    .X(\heichips25_can_lehmann_fsm/net844 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold846  (.A(\heichips25_can_lehmann_fsm/_0225_ ),
    .X(\heichips25_can_lehmann_fsm/net845 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold847  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[141] ),
    .X(\heichips25_can_lehmann_fsm/net846 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold848  (.A(\heichips25_can_lehmann_fsm/_0201_ ),
    .X(\heichips25_can_lehmann_fsm/net847 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold849  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[3] ),
    .X(\heichips25_can_lehmann_fsm/net848 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold850  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[188] ),
    .X(\heichips25_can_lehmann_fsm/net849 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold851  (.A(\heichips25_can_lehmann_fsm/_0248_ ),
    .X(\heichips25_can_lehmann_fsm/net850 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold852  (.A(\heichips25_can_lehmann_fsm/controller.const_data[9] ),
    .X(\heichips25_can_lehmann_fsm/net851 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold853  (.A(\heichips25_can_lehmann_fsm/_0069_ ),
    .X(\heichips25_can_lehmann_fsm/net852 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold854  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[181] ),
    .X(\heichips25_can_lehmann_fsm/net853 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold855  (.A(\heichips25_can_lehmann_fsm/_0241_ ),
    .X(\heichips25_can_lehmann_fsm/net854 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold856  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[163] ),
    .X(\heichips25_can_lehmann_fsm/net855 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold857  (.A(\heichips25_can_lehmann_fsm/_0223_ ),
    .X(\heichips25_can_lehmann_fsm/net856 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold858  (.A(\heichips25_can_lehmann_fsm/controller.const_data[16] ),
    .X(\heichips25_can_lehmann_fsm/net857 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold859  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[95] ),
    .X(\heichips25_can_lehmann_fsm/net858 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold860  (.A(\heichips25_can_lehmann_fsm/_0154_ ),
    .X(\heichips25_can_lehmann_fsm/net859 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold861  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[164] ),
    .X(\heichips25_can_lehmann_fsm/net860 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold862  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[81] ),
    .X(\heichips25_can_lehmann_fsm/net861 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold863  (.A(\heichips25_can_lehmann_fsm/_0141_ ),
    .X(\heichips25_can_lehmann_fsm/net862 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold864  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[99] ),
    .X(\heichips25_can_lehmann_fsm/net863 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold865  (.A(\heichips25_can_lehmann_fsm/_0159_ ),
    .X(\heichips25_can_lehmann_fsm/net864 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold866  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[61] ),
    .X(\heichips25_can_lehmann_fsm/net865 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold867  (.A(\heichips25_can_lehmann_fsm/_0120_ ),
    .X(\heichips25_can_lehmann_fsm/net866 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold868  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[175] ),
    .X(\heichips25_can_lehmann_fsm/net867 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold869  (.A(\heichips25_can_lehmann_fsm/_0234_ ),
    .X(\heichips25_can_lehmann_fsm/net868 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold870  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[80] ),
    .X(\heichips25_can_lehmann_fsm/net869 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold871  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[55] ),
    .X(\heichips25_can_lehmann_fsm/net870 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold872  (.A(\heichips25_can_lehmann_fsm/_0114_ ),
    .X(\heichips25_can_lehmann_fsm/net871 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold873  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[145] ),
    .X(\heichips25_can_lehmann_fsm/net872 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold874  (.A(\heichips25_can_lehmann_fsm/_0205_ ),
    .X(\heichips25_can_lehmann_fsm/net873 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold875  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[131] ),
    .X(\heichips25_can_lehmann_fsm/net874 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold876  (.A(\heichips25_can_lehmann_fsm/_0190_ ),
    .X(\heichips25_can_lehmann_fsm/net875 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold877  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[62] ),
    .X(\heichips25_can_lehmann_fsm/net876 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold878  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[8] ),
    .X(\heichips25_can_lehmann_fsm/net877 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold879  (.A(\heichips25_can_lehmann_fsm/_0268_ ),
    .X(\heichips25_can_lehmann_fsm/net878 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold880  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[48] ),
    .X(\heichips25_can_lehmann_fsm/net879 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold881  (.A(\heichips25_can_lehmann_fsm/_0108_ ),
    .X(\heichips25_can_lehmann_fsm/net880 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold882  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[177] ),
    .X(\heichips25_can_lehmann_fsm/net881 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold883  (.A(\heichips25_can_lehmann_fsm/_0236_ ),
    .X(\heichips25_can_lehmann_fsm/net882 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold884  (.A(\heichips25_can_lehmann_fsm/controller.const_data[31] ),
    .X(\heichips25_can_lehmann_fsm/net883 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold885  (.A(\heichips25_can_lehmann_fsm/_0090_ ),
    .X(\heichips25_can_lehmann_fsm/net884 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold886  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[133] ),
    .X(\heichips25_can_lehmann_fsm/net885 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold887  (.A(\heichips25_can_lehmann_fsm/_0192_ ),
    .X(\heichips25_can_lehmann_fsm/net886 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold888  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[135] ),
    .X(\heichips25_can_lehmann_fsm/net887 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold889  (.A(\heichips25_can_lehmann_fsm/_0195_ ),
    .X(\heichips25_can_lehmann_fsm/net888 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold890  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[153] ),
    .X(\heichips25_can_lehmann_fsm/net889 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold891  (.A(\heichips25_can_lehmann_fsm/_0212_ ),
    .X(\heichips25_can_lehmann_fsm/net890 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold892  (.A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[4] ),
    .X(\heichips25_sap3/net891 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold893  (.A(\heichips25_sap3/_0177_ ),
    .X(\heichips25_sap3/net892 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold894  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[89] ),
    .X(\heichips25_can_lehmann_fsm/net893 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold895  (.A(\heichips25_can_lehmann_fsm/_0149_ ),
    .X(\heichips25_can_lehmann_fsm/net894 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold896  (.A(\heichips25_can_lehmann_fsm/controller.const_data[3] ),
    .X(\heichips25_can_lehmann_fsm/net895 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold897  (.A(\heichips25_can_lehmann_fsm/_0062_ ),
    .X(\heichips25_can_lehmann_fsm/net896 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold898  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[144] ),
    .X(\heichips25_can_lehmann_fsm/net897 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold899  (.A(\heichips25_can_lehmann_fsm/controller.const_data[19] ),
    .X(\heichips25_can_lehmann_fsm/net898 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold900  (.A(\heichips25_can_lehmann_fsm/_0079_ ),
    .X(\heichips25_can_lehmann_fsm/net899 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold901  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[73] ),
    .X(\heichips25_can_lehmann_fsm/net900 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold902  (.A(\heichips25_can_lehmann_fsm/_0132_ ),
    .X(\heichips25_can_lehmann_fsm/net901 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold903  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[132] ),
    .X(\heichips25_can_lehmann_fsm/net902 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold904  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[74] ),
    .X(\heichips25_can_lehmann_fsm/net903 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold905  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[111] ),
    .X(\heichips25_can_lehmann_fsm/net904 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold906  (.A(\heichips25_can_lehmann_fsm/_0171_ ),
    .X(\heichips25_can_lehmann_fsm/net905 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold907  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[169] ),
    .X(\heichips25_can_lehmann_fsm/net906 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold908  (.A(\heichips25_can_lehmann_fsm/_0228_ ),
    .X(\heichips25_can_lehmann_fsm/net907 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold909  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[7] ),
    .X(\heichips25_can_lehmann_fsm/net908 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold910  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[75] ),
    .X(\heichips25_can_lehmann_fsm/net909 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold911  (.A(\heichips25_can_lehmann_fsm/_0135_ ),
    .X(\heichips25_can_lehmann_fsm/net910 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold912  (.A(\heichips25_can_lehmann_fsm/controller.const_data[18] ),
    .X(\heichips25_can_lehmann_fsm/net911 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold913  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[32] ),
    .X(\heichips25_can_lehmann_fsm/net912 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold914  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[63] ),
    .X(\heichips25_can_lehmann_fsm/net913 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold915  (.A(\heichips25_can_lehmann_fsm/_0123_ ),
    .X(\heichips25_can_lehmann_fsm/net914 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold916  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[176] ),
    .X(\heichips25_can_lehmann_fsm/net915 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold917  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[51] ),
    .X(\heichips25_can_lehmann_fsm/net916 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold918  (.A(\heichips25_can_lehmann_fsm/_0111_ ),
    .X(\heichips25_can_lehmann_fsm/net917 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold919  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[157] ),
    .X(\heichips25_can_lehmann_fsm/net918 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold920  (.A(\heichips25_can_lehmann_fsm/_0216_ ),
    .X(\heichips25_can_lehmann_fsm/net919 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold921  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[170] ),
    .X(\heichips25_can_lehmann_fsm/net920 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold922  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[134] ),
    .X(\heichips25_can_lehmann_fsm/net921 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold923  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[33] ),
    .X(\heichips25_can_lehmann_fsm/net922 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold924  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[178] ),
    .X(\heichips25_can_lehmann_fsm/net923 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold925  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[180] ),
    .X(\heichips25_can_lehmann_fsm/net924 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold926  (.A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[3] ),
    .X(\heichips25_sap3/net925 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold927  (.A(\heichips25_sap3/_0176_ ),
    .X(\heichips25_sap3/net926 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold928  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[143] ),
    .X(\heichips25_can_lehmann_fsm/net927 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold929  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[161] ),
    .X(\heichips25_can_lehmann_fsm/net928 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold930  (.A(\heichips25_can_lehmann_fsm/_0220_ ),
    .X(\heichips25_can_lehmann_fsm/net929 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold931  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[142] ),
    .X(\heichips25_can_lehmann_fsm/net930 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold932  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[171] ),
    .X(\heichips25_can_lehmann_fsm/net931 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold933  (.A(\heichips25_can_lehmann_fsm/_0231_ ),
    .X(\heichips25_can_lehmann_fsm/net932 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold934  (.A(\heichips25_can_lehmann_fsm/controller.const_data[4] ),
    .X(\heichips25_can_lehmann_fsm/net933 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold935  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[113] ),
    .X(\heichips25_can_lehmann_fsm/net934 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold936  (.A(\heichips25_can_lehmann_fsm/_0172_ ),
    .X(\heichips25_can_lehmann_fsm/net935 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold937  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[96] ),
    .X(\heichips25_can_lehmann_fsm/net936 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold938  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[87] ),
    .X(\heichips25_can_lehmann_fsm/net937 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold939  (.A(\heichips25_can_lehmann_fsm/_0146_ ),
    .X(\heichips25_can_lehmann_fsm/net938 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold940  (.A(\heichips25_can_lehmann_fsm/controller.const_data[21] ),
    .X(\heichips25_can_lehmann_fsm/net939 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold941  (.A(\heichips25_can_lehmann_fsm/_0080_ ),
    .X(\heichips25_can_lehmann_fsm/net940 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold942  (.A(\heichips25_can_lehmann_fsm/controller.const_data[22] ),
    .X(\heichips25_can_lehmann_fsm/net941 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold943  (.A(\heichips25_can_lehmann_fsm/controller.const_data[25] ),
    .X(\heichips25_can_lehmann_fsm/net942 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold944  (.A(\heichips25_can_lehmann_fsm/_0084_ ),
    .X(\heichips25_can_lehmann_fsm/net943 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold945  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[6] ),
    .X(\heichips25_can_lehmann_fsm/net944 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold946  (.A(\heichips25_can_lehmann_fsm/_0265_ ),
    .X(\heichips25_can_lehmann_fsm/net945 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold947  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[137] ),
    .X(\heichips25_can_lehmann_fsm/net946 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold948  (.A(\heichips25_can_lehmann_fsm/_0196_ ),
    .X(\heichips25_can_lehmann_fsm/net947 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold949  (.A(\heichips25_can_lehmann_fsm/controller.const_data[27] ),
    .X(\heichips25_can_lehmann_fsm/net948 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold950  (.A(\heichips25_can_lehmann_fsm/_0086_ ),
    .X(\heichips25_can_lehmann_fsm/net949 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold951  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[98] ),
    .X(\heichips25_can_lehmann_fsm/net950 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold952  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[196] ),
    .X(\heichips25_can_lehmann_fsm/net951 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold953  (.A(\heichips25_can_lehmann_fsm/_0256_ ),
    .X(\heichips25_can_lehmann_fsm/net952 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold954  (.A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[6] ),
    .X(\heichips25_sap3/net953 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold955  (.A(\heichips25_sap3/_0179_ ),
    .X(\heichips25_sap3/net954 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold956  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[57] ),
    .X(\heichips25_can_lehmann_fsm/net955 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold957  (.A(\heichips25_can_lehmann_fsm/_0116_ ),
    .X(\heichips25_can_lehmann_fsm/net956 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold958  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[139] ),
    .X(\heichips25_can_lehmann_fsm/net957 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold959  (.A(\heichips25_can_lehmann_fsm/_0199_ ),
    .X(\heichips25_can_lehmann_fsm/net958 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold960  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[140] ),
    .X(\heichips25_can_lehmann_fsm/net959 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold961  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[192] ),
    .X(\heichips25_can_lehmann_fsm/net960 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold962  (.A(\heichips25_can_lehmann_fsm/_0252_ ),
    .X(\heichips25_can_lehmann_fsm/net961 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold963  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[88] ),
    .X(\heichips25_can_lehmann_fsm/net962 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold964  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[154] ),
    .X(\heichips25_can_lehmann_fsm/net963 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold965  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[158] ),
    .X(\heichips25_can_lehmann_fsm/net964 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold966  (.A(\heichips25_can_lehmann_fsm/controller.const_data[23] ),
    .X(\heichips25_can_lehmann_fsm/net965 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold967  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[77] ),
    .X(\heichips25_can_lehmann_fsm/net966 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold968  (.A(\heichips25_can_lehmann_fsm/_0136_ ),
    .X(\heichips25_can_lehmann_fsm/net967 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold969  (.A(\heichips25_can_lehmann_fsm/controller.const_data[24] ),
    .X(\heichips25_can_lehmann_fsm/net968 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold970  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[110] ),
    .X(\heichips25_can_lehmann_fsm/net969 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold971  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[107] ),
    .X(\heichips25_can_lehmann_fsm/net970 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold972  (.A(\heichips25_can_lehmann_fsm/_0167_ ),
    .X(\heichips25_can_lehmann_fsm/net971 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold973  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[138] ),
    .X(\heichips25_can_lehmann_fsm/net972 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold974  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[56] ),
    .X(\heichips25_can_lehmann_fsm/net973 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold975  (.A(\heichips25_can_lehmann_fsm/controller.const_data[8] ),
    .X(\heichips25_can_lehmann_fsm/net974 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold976  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[78] ),
    .X(\heichips25_can_lehmann_fsm/net975 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold977  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[50] ),
    .X(\heichips25_can_lehmann_fsm/net976 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold978  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[49] ),
    .X(\heichips25_can_lehmann_fsm/net977 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold979  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[151] ),
    .X(\heichips25_can_lehmann_fsm/net978 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold980  (.A(\heichips25_can_lehmann_fsm/_0211_ ),
    .X(\heichips25_can_lehmann_fsm/net979 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold981  (.A(\heichips25_can_lehmann_fsm/controller.const_data[26] ),
    .X(\heichips25_can_lehmann_fsm/net980 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold982  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[85] ),
    .X(\heichips25_can_lehmann_fsm/net981 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold983  (.A(\heichips25_can_lehmann_fsm/_0145_ ),
    .X(\heichips25_can_lehmann_fsm/net982 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold984  (.A(\heichips25_can_lehmann_fsm/controller.const_data[28] ),
    .X(\heichips25_can_lehmann_fsm/net983 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold985  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[150] ),
    .X(\heichips25_can_lehmann_fsm/net984 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold986  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[149] ),
    .X(\heichips25_can_lehmann_fsm/net985 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold987  (.A(\heichips25_can_lehmann_fsm/_0208_ ),
    .X(\heichips25_can_lehmann_fsm/net986 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold988  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[35] ),
    .X(\heichips25_can_lehmann_fsm/net987 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold989  (.A(\heichips25_can_lehmann_fsm/_0094_ ),
    .X(\heichips25_can_lehmann_fsm/net988 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold990  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[58] ),
    .X(\heichips25_can_lehmann_fsm/net989 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold991  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[185] ),
    .X(\heichips25_can_lehmann_fsm/net990 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold992  (.A(\heichips25_can_lehmann_fsm/_0244_ ),
    .X(\heichips25_can_lehmann_fsm/net991 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold993  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[97] ),
    .X(\heichips25_can_lehmann_fsm/net992 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold994  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[198] ),
    .X(\heichips25_can_lehmann_fsm/net993 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold995  (.A(\heichips25_can_lehmann_fsm/_0258_ ),
    .X(\heichips25_can_lehmann_fsm/net994 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold996  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[159] ),
    .X(\heichips25_can_lehmann_fsm/net995 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold997  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[69] ),
    .X(\heichips25_can_lehmann_fsm/net996 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold998  (.A(\heichips25_can_lehmann_fsm/_0129_ ),
    .X(\heichips25_can_lehmann_fsm/net997 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold999  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[183] ),
    .X(\heichips25_can_lehmann_fsm/net998 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1000  (.A(\heichips25_can_lehmann_fsm/_0242_ ),
    .X(\heichips25_can_lehmann_fsm/net999 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1001  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[45] ),
    .X(\heichips25_can_lehmann_fsm/net1000 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1002  (.A(\heichips25_can_lehmann_fsm/_0105_ ),
    .X(\heichips25_can_lehmann_fsm/net1001 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1003  (.A(\heichips25_can_lehmann_fsm/controller.const_data[15] ),
    .X(\heichips25_can_lehmann_fsm/net1002 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1004  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[53] ),
    .X(\heichips25_can_lehmann_fsm/net1003 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1005  (.A(\heichips25_can_lehmann_fsm/_0113_ ),
    .X(\heichips25_can_lehmann_fsm/net1004 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1006  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[106] ),
    .X(\heichips25_can_lehmann_fsm/net1005 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1007  (.A(\heichips25_can_lehmann_fsm/controller.const_data[11] ),
    .X(\heichips25_can_lehmann_fsm/net1006 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1008  (.A(\heichips25_can_lehmann_fsm/_0070_ ),
    .X(\heichips25_can_lehmann_fsm/net1007 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1009  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[67] ),
    .X(\heichips25_can_lehmann_fsm/net1008 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1010  (.A(\heichips25_can_lehmann_fsm/_0126_ ),
    .X(\heichips25_can_lehmann_fsm/net1009 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1011  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[160] ),
    .X(\heichips25_can_lehmann_fsm/net1010 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold1012  (.A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[5] ),
    .X(\heichips25_sap3/net1011 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold1013  (.A(\heichips25_sap3/_0178_ ),
    .X(\heichips25_sap3/net1012 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1014  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[103] ),
    .X(\heichips25_can_lehmann_fsm/net1013 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1015  (.A(\heichips25_can_lehmann_fsm/_0163_ ),
    .X(\heichips25_can_lehmann_fsm/net1014 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1016  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[40] ),
    .X(\heichips25_can_lehmann_fsm/net1015 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1017  (.A(\heichips25_can_lehmann_fsm/_0100_ ),
    .X(\heichips25_can_lehmann_fsm/net1016 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1018  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[127] ),
    .X(\heichips25_can_lehmann_fsm/net1017 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1019  (.A(\heichips25_can_lehmann_fsm/_0186_ ),
    .X(\heichips25_can_lehmann_fsm/net1018 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold1020  (.A(\heichips25_sap3/u_ser.bit_pos[2] ),
    .X(\heichips25_sap3/net1019 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold1021  (.A(\heichips25_sap3/_0017_ ),
    .X(\heichips25_sap3/net1020 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1022  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[155] ),
    .X(\heichips25_can_lehmann_fsm/net1021 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1023  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[147] ),
    .X(\heichips25_can_lehmann_fsm/net1022 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1024  (.A(\heichips25_can_lehmann_fsm/_0206_ ),
    .X(\heichips25_can_lehmann_fsm/net1023 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1025  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[68] ),
    .X(\heichips25_can_lehmann_fsm/net1024 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1026  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[109] ),
    .X(\heichips25_can_lehmann_fsm/net1025 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1027  (.A(\heichips25_can_lehmann_fsm/_0168_ ),
    .X(\heichips25_can_lehmann_fsm/net1026 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1028  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[121] ),
    .X(\heichips25_can_lehmann_fsm/net1027 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1029  (.A(\heichips25_can_lehmann_fsm/_0180_ ),
    .X(\heichips25_can_lehmann_fsm/net1028 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1030  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[195] ),
    .X(\heichips25_can_lehmann_fsm/net1029 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1031  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[148] ),
    .X(\heichips25_can_lehmann_fsm/net1030 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold1032  (.A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[7] ),
    .X(\heichips25_sap3/net1031 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold1033  (.A(\heichips25_sap3/_0180_ ),
    .X(\heichips25_sap3/net1032 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1034  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[184] ),
    .X(\heichips25_can_lehmann_fsm/net1033 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1035  (.A(\heichips25_can_lehmann_fsm/controller.const_data[12] ),
    .X(\heichips25_can_lehmann_fsm/net1034 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1036  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[123] ),
    .X(\heichips25_can_lehmann_fsm/net1035 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1037  (.A(\heichips25_can_lehmann_fsm/_0182_ ),
    .X(\heichips25_can_lehmann_fsm/net1036 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1038  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[114] ),
    .X(\heichips25_can_lehmann_fsm/net1037 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1039  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[128] ),
    .X(\heichips25_can_lehmann_fsm/net1038 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1040  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[197] ),
    .X(\heichips25_can_lehmann_fsm/net1039 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1041  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[122] ),
    .X(\heichips25_can_lehmann_fsm/net1040 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1042  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[71] ),
    .X(\heichips25_can_lehmann_fsm/net1041 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1043  (.A(\heichips25_can_lehmann_fsm/_0130_ ),
    .X(\heichips25_can_lehmann_fsm/net1042 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1044  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[21] ),
    .X(\heichips25_can_lehmann_fsm/net1043 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1045  (.A(\heichips25_can_lehmann_fsm/_0280_ ),
    .X(\heichips25_can_lehmann_fsm/net1044 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1046  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[125] ),
    .X(\heichips25_can_lehmann_fsm/net1045 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1047  (.A(\heichips25_can_lehmann_fsm/_0185_ ),
    .X(\heichips25_can_lehmann_fsm/net1046 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1048  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[91] ),
    .X(\heichips25_can_lehmann_fsm/net1047 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1049  (.A(\heichips25_can_lehmann_fsm/_0151_ ),
    .X(\heichips25_can_lehmann_fsm/net1048 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1050  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[79] ),
    .X(\heichips25_can_lehmann_fsm/net1049 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1051  (.A(\heichips25_can_lehmann_fsm/controller.const_data[13] ),
    .X(\heichips25_can_lehmann_fsm/net1050 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1052  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[19] ),
    .X(\heichips25_can_lehmann_fsm/net1051 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1053  (.A(\heichips25_can_lehmann_fsm/_0278_ ),
    .X(\heichips25_can_lehmann_fsm/net1052 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1054  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[156] ),
    .X(\heichips25_can_lehmann_fsm/net1053 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1055  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[90] ),
    .X(\heichips25_can_lehmann_fsm/net1054 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1056  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[44] ),
    .X(\heichips25_can_lehmann_fsm/net1055 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1057  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[65] ),
    .X(\heichips25_can_lehmann_fsm/net1056 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1058  (.A(\heichips25_can_lehmann_fsm/_0124_ ),
    .X(\heichips25_can_lehmann_fsm/net1057 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold1059  (.A(\heichips25_sap3/regFile_serial ),
    .X(\heichips25_sap3/net1058 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold1060  (.A(\heichips25_sap3/_0168_ ),
    .X(\heichips25_sap3/net1059 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1061  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[115] ),
    .X(\heichips25_can_lehmann_fsm/net1060 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1062  (.A(\heichips25_can_lehmann_fsm/_0175_ ),
    .X(\heichips25_can_lehmann_fsm/net1061 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1063  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[93] ),
    .X(\heichips25_can_lehmann_fsm/net1062 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1064  (.A(\heichips25_can_lehmann_fsm/_0153_ ),
    .X(\heichips25_can_lehmann_fsm/net1063 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold1065  (.A(\heichips25_sap3/u_ser.state[1] ),
    .X(\heichips25_sap3/net1064 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold1066  (.A(\heichips25_sap3/_0287_ ),
    .X(\heichips25_sap3/net1065 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1067  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[38] ),
    .X(\heichips25_can_lehmann_fsm/net1066 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1068  (.A(\heichips25_can_lehmann_fsm/_0098_ ),
    .X(\heichips25_can_lehmann_fsm/net1067 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1069  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[34] ),
    .X(\heichips25_can_lehmann_fsm/net1068 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1070  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[66] ),
    .X(\heichips25_can_lehmann_fsm/net1069 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1071  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[84] ),
    .X(\heichips25_can_lehmann_fsm/net1070 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold1072  (.A(\heichips25_sap3/u_ser.bit_pos[0] ),
    .X(\heichips25_sap3/net1071 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold1073  (.A(\heichips25_sap3/_1356_ ),
    .X(\heichips25_sap3/net1072 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold1074  (.A(\heichips25_sap3/_0188_ ),
    .X(\heichips25_sap3/net1073 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1075  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[190] ),
    .X(\heichips25_can_lehmann_fsm/net1074 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1076  (.A(\heichips25_can_lehmann_fsm/_0250_ ),
    .X(\heichips25_can_lehmann_fsm/net1075 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1077  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[191] ),
    .X(\heichips25_can_lehmann_fsm/net1076 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1078  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[117] ),
    .X(\heichips25_can_lehmann_fsm/net1077 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1079  (.A(\heichips25_can_lehmann_fsm/_0176_ ),
    .X(\heichips25_can_lehmann_fsm/net1078 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1080  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[102] ),
    .X(\heichips25_can_lehmann_fsm/net1079 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1081  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[39] ),
    .X(\heichips25_can_lehmann_fsm/net1080 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1082  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[36] ),
    .X(\heichips25_can_lehmann_fsm/net1081 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1083  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[118] ),
    .X(\heichips25_can_lehmann_fsm/net1082 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1084  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[129] ),
    .X(\heichips25_can_lehmann_fsm/net1083 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1085  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[20] ),
    .X(\heichips25_can_lehmann_fsm/net1084 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1086  (.A(\heichips25_can_lehmann_fsm/controller.const_data[29] ),
    .X(\heichips25_can_lehmann_fsm/net1085 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1087  (.A(\heichips25_can_lehmann_fsm/_0089_ ),
    .X(\heichips25_can_lehmann_fsm/net1086 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1088  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[186] ),
    .X(\heichips25_can_lehmann_fsm/net1087 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1089  (.A(\heichips25_can_lehmann_fsm/controller.const_data[7] ),
    .X(\heichips25_can_lehmann_fsm/net1088 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1090  (.A(\heichips25_can_lehmann_fsm/_0066_ ),
    .X(\heichips25_can_lehmann_fsm/net1089 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1091  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[162] ),
    .X(\heichips25_can_lehmann_fsm/net1090 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1092  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[130] ),
    .X(\heichips25_can_lehmann_fsm/net1091 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1093  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[92] ),
    .X(\heichips25_can_lehmann_fsm/net1092 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1094  (.A(\heichips25_can_lehmann_fsm/controller.const_data[1] ),
    .X(\heichips25_can_lehmann_fsm/net1093 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1095  (.A(\heichips25_can_lehmann_fsm/_0060_ ),
    .X(\heichips25_can_lehmann_fsm/net1094 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1096  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[47] ),
    .X(\heichips25_can_lehmann_fsm/net1095 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1097  (.A(\heichips25_can_lehmann_fsm/_0106_ ),
    .X(\heichips25_can_lehmann_fsm/net1096 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1098  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[105] ),
    .X(\heichips25_can_lehmann_fsm/net1097 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1099  (.A(\heichips25_can_lehmann_fsm/_0164_ ),
    .X(\heichips25_can_lehmann_fsm/net1098 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1100  (.A(\heichips25_can_lehmann_fsm/controller.const_data[5] ),
    .X(\heichips25_can_lehmann_fsm/net1099 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1101  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[59] ),
    .X(\heichips25_can_lehmann_fsm/net1100 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1102  (.A(\heichips25_can_lehmann_fsm/_0119_ ),
    .X(\heichips25_can_lehmann_fsm/net1101 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1103  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[72] ),
    .X(\heichips25_can_lehmann_fsm/net1102 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1104  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[119] ),
    .X(\heichips25_can_lehmann_fsm/net1103 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1105  (.A(\heichips25_can_lehmann_fsm/_0179_ ),
    .X(\heichips25_can_lehmann_fsm/net1104 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold1106  (.A(\heichips25_sap3/u_ser.shadow_reg[6] ),
    .X(\heichips25_sap3/net1105 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1107  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[101] ),
    .X(\heichips25_can_lehmann_fsm/net1106 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1108  (.A(\heichips25_can_lehmann_fsm/_0160_ ),
    .X(\heichips25_can_lehmann_fsm/net1107 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1109  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[83] ),
    .X(\heichips25_can_lehmann_fsm/net1108 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1110  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[124] ),
    .X(\heichips25_can_lehmann_fsm/net1109 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1111  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[42] ),
    .X(\heichips25_can_lehmann_fsm/net1110 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1112  (.A(\heichips25_can_lehmann_fsm/_0101_ ),
    .X(\heichips25_can_lehmann_fsm/net1111 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold1113  (.A(\heichips25_sap3/u_ser.shadow_reg[7] ),
    .X(\heichips25_sap3/net1112 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1114  (.A(\heichips25_can_lehmann_fsm/controller.const_data[6] ),
    .X(\heichips25_can_lehmann_fsm/net1113 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1115  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[189] ),
    .X(\heichips25_can_lehmann_fsm/net1114 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1116  (.A(\heichips25_can_lehmann_fsm/controller.const_data[14] ),
    .X(\heichips25_can_lehmann_fsm/net1115 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1117  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[22] ),
    .X(\heichips25_can_lehmann_fsm/net1116 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1118  (.A(\heichips25_can_lehmann_fsm/controller.extended_then_action[3] ),
    .X(\heichips25_can_lehmann_fsm/net1117 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1119  (.A(\heichips25_can_lehmann_fsm/_0275_ ),
    .X(\heichips25_can_lehmann_fsm/net1118 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold1120  (.A(\heichips25_sap3/u_ser.shadow_reg[3] ),
    .X(\heichips25_sap3/net1119 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold1121  (.A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[2] ),
    .X(\heichips25_sap3/net1120 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold1122  (.A(\heichips25_sap3/u_ser.shadow_reg[1] ),
    .X(\heichips25_sap3/net1121 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1123  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[167] ),
    .X(\heichips25_can_lehmann_fsm/net1122 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1124  (.A(\heichips25_can_lehmann_fsm/_0226_ ),
    .X(\heichips25_can_lehmann_fsm/net1123 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold1125  (.A(\heichips25_sap3/u_ser.shadow_reg[5] ),
    .X(\heichips25_sap3/net1124 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold1126  (.A(\heichips25_sap3/_0195_ ),
    .X(\heichips25_sap3/net1125 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1127  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[43] ),
    .X(\heichips25_can_lehmann_fsm/net1126 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1128  (.A(\heichips25_can_lehmann_fsm/controller.extended_then_action[2] ),
    .X(\heichips25_can_lehmann_fsm/net1127 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold1129  (.A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[0] ),
    .X(\heichips25_sap3/net1128 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1130  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[179] ),
    .X(\heichips25_can_lehmann_fsm/net1129 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold1131  (.A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.state[1] ),
    .X(\heichips25_sap3/net1130 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold1132  (.A(\heichips25_sap3/_0291_ ),
    .X(\heichips25_sap3/net1131 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1133  (.A(\heichips25_can_lehmann_fsm/controller.extended_state[1] ),
    .X(\heichips25_can_lehmann_fsm/net1132 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1134  (.A(\heichips25_can_lehmann_fsm/_0284_ ),
    .X(\heichips25_can_lehmann_fsm/net1133 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1135  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[168] ),
    .X(\heichips25_can_lehmann_fsm/net1134 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1136  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[82] ),
    .X(\heichips25_can_lehmann_fsm/net1135 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1137  (.A(\heichips25_can_lehmann_fsm/controller.const_data[2] ),
    .X(\heichips25_can_lehmann_fsm/net1136 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1138  (.A(\heichips25_can_lehmann_fsm/controller.extended_state[2] ),
    .X(\heichips25_can_lehmann_fsm/net1137 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold1139  (.A(\heichips25_sap3/u_ser.bit_pos[1] ),
    .X(\heichips25_sap3/net1138 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1140  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[173] ),
    .X(\heichips25_can_lehmann_fsm/net1139 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1141  (.A(\heichips25_can_lehmann_fsm/_0232_ ),
    .X(\heichips25_can_lehmann_fsm/net1140 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold1142  (.A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[1] ),
    .X(\heichips25_sap3/net1141 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1143  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.extended_word[23] ),
    .X(\heichips25_can_lehmann_fsm/net1142 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold1144  (.A(\heichips25_sap3/u_ser.shadow_reg[4] ),
    .X(\heichips25_sap3/net1143 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold1145  (.A(\heichips25_sap3/_0194_ ),
    .X(\heichips25_sap3/net1144 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold1146  (.A(\heichips25_sap3/u_ser.shadow_reg[0] ),
    .X(\heichips25_sap3/net1145 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1147  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[187] ),
    .X(\heichips25_can_lehmann_fsm/net1146 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1148  (.A(\heichips25_can_lehmann_fsm/controller.extended_then_action[1] ),
    .X(\heichips25_can_lehmann_fsm/net1147 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1149  (.A(\heichips25_can_lehmann_fsm/controller.extended_state[0] ),
    .X(\heichips25_can_lehmann_fsm/net1148 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold1150  (.A(\heichips25_sap3/u_ser.shadow_reg[2] ),
    .X(\heichips25_sap3/net1149 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1151  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[174] ),
    .X(\heichips25_can_lehmann_fsm/net1150 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1152  (.A(\heichips25_can_lehmann_fsm/controller.extended_then_action[0] ),
    .X(\heichips25_can_lehmann_fsm/net1151 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1153  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[194] ),
    .X(\heichips25_can_lehmann_fsm/net1152 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1154  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[193] ),
    .X(\heichips25_can_lehmann_fsm/net1153 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1155  (.A(\heichips25_can_lehmann_fsm/controller.extended_cond.opcode[2] ),
    .X(\heichips25_can_lehmann_fsm/net1154 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1156  (.A(\heichips25_can_lehmann_fsm/controller.extended_then_action[5] ),
    .X(\heichips25_can_lehmann_fsm/net1155 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1157  (.A(\heichips25_can_lehmann_fsm/_0277_ ),
    .X(\heichips25_can_lehmann_fsm/net1156 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1158  (.A(\heichips25_can_lehmann_fsm/controller.extended_then_action[4] ),
    .X(\heichips25_can_lehmann_fsm/net1157 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1159  (.A(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[13] ),
    .X(\heichips25_can_lehmann_fsm/net1158 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1160  (.A(\heichips25_can_lehmann_fsm/_0056_ ),
    .X(\heichips25_can_lehmann_fsm/net1159 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1161  (.A(\heichips25_can_lehmann_fsm/controller.extended_jump_target[0] ),
    .X(\heichips25_can_lehmann_fsm/net1160 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1162  (.A(\heichips25_can_lehmann_fsm/_0259_ ),
    .X(\heichips25_can_lehmann_fsm/net1161 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold1163  (.A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos[1] ),
    .X(\heichips25_sap3/net1162 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold1164  (.A(\heichips25_sap3/_1255_ ),
    .X(\heichips25_sap3/net1163 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1165  (.A(\heichips25_can_lehmann_fsm/controller.extended_jump_target[2] ),
    .X(\heichips25_can_lehmann_fsm/net1164 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1166  (.A(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[11] ),
    .X(\heichips25_can_lehmann_fsm/net1165 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1167  (.A(\heichips25_can_lehmann_fsm/_0054_ ),
    .X(\heichips25_can_lehmann_fsm/net1166 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1168  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[37] ),
    .X(\heichips25_can_lehmann_fsm/net1167 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1169  (.A(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[15] ),
    .X(\heichips25_can_lehmann_fsm/net1168 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1170  (.A(\heichips25_can_lehmann_fsm/_0621_ ),
    .X(\heichips25_can_lehmann_fsm/net1169 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1171  (.A(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[9] ),
    .X(\heichips25_can_lehmann_fsm/net1170 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1172  (.A(\heichips25_can_lehmann_fsm/_0052_ ),
    .X(\heichips25_can_lehmann_fsm/net1171 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1173  (.A(\heichips25_can_lehmann_fsm/controller.extended_jump_target[1] ),
    .X(\heichips25_can_lehmann_fsm/net1172 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1174  (.A(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[3] ),
    .X(\heichips25_can_lehmann_fsm/net1173 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1175  (.A(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[1] ),
    .X(\heichips25_can_lehmann_fsm/net1174 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1176  (.A(\heichips25_can_lehmann_fsm/_0044_ ),
    .X(\heichips25_can_lehmann_fsm/net1175 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold1177  (.A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos[0] ),
    .X(\heichips25_sap3/net1176 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1178  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[52] ),
    .X(\heichips25_can_lehmann_fsm/net1177 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold1179  (.A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.word_index[1] ),
    .X(\heichips25_sap3/net1178 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold1180  (.A(\heichips25_sap3/_0182_ ),
    .X(\heichips25_sap3/net1179 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1181  (.A(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[9] ),
    .X(\heichips25_can_lehmann_fsm/net1180 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1182  (.A(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[5] ),
    .X(\heichips25_can_lehmann_fsm/net1181 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1183  (.A(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[7] ),
    .X(\heichips25_can_lehmann_fsm/net1182 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1184  (.A(\heichips25_can_lehmann_fsm/controller.const_data[20] ),
    .X(\heichips25_can_lehmann_fsm/net1183 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1185  (.A(\heichips25_can_lehmann_fsm/_0576_ ),
    .X(\heichips25_can_lehmann_fsm/net1184 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1186  (.A(\heichips25_can_lehmann_fsm/_0047_ ),
    .X(\heichips25_can_lehmann_fsm/net1185 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1187  (.A(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[11] ),
    .X(\heichips25_can_lehmann_fsm/net1186 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1188  (.A(\heichips25_can_lehmann_fsm/_0038_ ),
    .X(\heichips25_can_lehmann_fsm/net1187 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1189  (.A(\heichips25_can_lehmann_fsm/controller.const_data[30] ),
    .X(\heichips25_can_lehmann_fsm/net1188 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1190  (.A(\heichips25_can_lehmann_fsm/_0618_ ),
    .X(\heichips25_can_lehmann_fsm/net1189 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1191  (.A(\heichips25_can_lehmann_fsm/_0057_ ),
    .X(\heichips25_can_lehmann_fsm/net1190 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1192  (.A(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[8] ),
    .X(\heichips25_can_lehmann_fsm/net1191 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1193  (.A(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[6] ),
    .X(\heichips25_can_lehmann_fsm/net1192 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1194  (.A(\heichips25_can_lehmann_fsm/_0033_ ),
    .X(\heichips25_can_lehmann_fsm/net1193 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1195  (.A(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[6] ),
    .X(\heichips25_can_lehmann_fsm/net1194 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1196  (.A(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[2] ),
    .X(\heichips25_can_lehmann_fsm/net1195 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1197  (.A(\heichips25_can_lehmann_fsm/_0045_ ),
    .X(\heichips25_can_lehmann_fsm/net1196 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold1198  (.A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.word_index[0] ),
    .X(\heichips25_sap3/net1197 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1199  (.A(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[7] ),
    .X(\heichips25_can_lehmann_fsm/net1198 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1200  (.A(\heichips25_can_lehmann_fsm/_0034_ ),
    .X(\heichips25_can_lehmann_fsm/net1199 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1201  (.A(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[12] ),
    .X(\heichips25_can_lehmann_fsm/net1200 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1202  (.A(\heichips25_can_lehmann_fsm/_0609_ ),
    .X(\heichips25_can_lehmann_fsm/net1201 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1203  (.A(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[3] ),
    .X(\heichips25_can_lehmann_fsm/net1202 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1204  (.A(\heichips25_can_lehmann_fsm/_0030_ ),
    .X(\heichips25_can_lehmann_fsm/net1203 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1205  (.A(\heichips25_can_lehmann_fsm/controller.const_data[0] ),
    .X(\heichips25_can_lehmann_fsm/net1204 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1206  (.A(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[15] ),
    .X(\heichips25_can_lehmann_fsm/net1205 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1207  (.A(\heichips25_can_lehmann_fsm/_0042_ ),
    .X(\heichips25_can_lehmann_fsm/net1206 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1208  (.A(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[10] ),
    .X(\heichips25_can_lehmann_fsm/net1207 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1209  (.A(\heichips25_can_lehmann_fsm/_0037_ ),
    .X(\heichips25_can_lehmann_fsm/net1208 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1210  (.A(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[10] ),
    .X(\heichips25_can_lehmann_fsm/net1209 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1211  (.A(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[5] ),
    .X(\heichips25_can_lehmann_fsm/net1210 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1212  (.A(\heichips25_can_lehmann_fsm/_0032_ ),
    .X(\heichips25_can_lehmann_fsm/net1211 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1213  (.A(\heichips25_can_lehmann_fsm/controller.counter2.counter_1[0] ),
    .X(\heichips25_can_lehmann_fsm/net1212 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1214  (.A(\heichips25_can_lehmann_fsm/controller.output_controller.keep[2] ),
    .X(\heichips25_can_lehmann_fsm/net1213 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1215  (.A(\heichips25_can_lehmann_fsm/_0288_ ),
    .X(\heichips25_can_lehmann_fsm/net1214 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1216  (.A(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[2] ),
    .X(\heichips25_can_lehmann_fsm/net1215 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1217  (.A(\heichips25_can_lehmann_fsm/_0029_ ),
    .X(\heichips25_can_lehmann_fsm/net1216 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1218  (.A(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[13] ),
    .X(\heichips25_can_lehmann_fsm/net1217 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1219  (.A(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[8] ),
    .X(\heichips25_can_lehmann_fsm/net1218 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1220  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[2] ),
    .X(\heichips25_can_lehmann_fsm/net1219 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1221  (.A(\heichips25_can_lehmann_fsm/_0022_ ),
    .X(\heichips25_can_lehmann_fsm/net1220 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1222  (.A(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[14] ),
    .X(\heichips25_can_lehmann_fsm/net1221 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1223  (.A(\heichips25_can_lehmann_fsm/_0041_ ),
    .X(\heichips25_can_lehmann_fsm/net1222 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold1224  (.A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.word_index[3] ),
    .X(\heichips25_sap3/net1223 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold1225  (.A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.word_index[2] ),
    .X(\heichips25_sap3/net1224 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold1226  (.A(\heichips25_sap3/u_ser.state[1] ),
    .X(\heichips25_sap3/net1225 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1227  (.A(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[0] ),
    .X(\heichips25_can_lehmann_fsm/net1226 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1228  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[23] ),
    .X(\heichips25_can_lehmann_fsm/net1227 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1229  (.A(\heichips25_can_lehmann_fsm/_0017_ ),
    .X(\heichips25_can_lehmann_fsm/net1228 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1230  (.A(\heichips25_can_lehmann_fsm/controller.extended_cond.opcode[1] ),
    .X(\heichips25_can_lehmann_fsm/net1229 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1231  (.A(\heichips25_can_lehmann_fsm/_0269_ ),
    .X(\heichips25_can_lehmann_fsm/net1230 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1232  (.A(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[12] ),
    .X(\heichips25_can_lehmann_fsm/net1231 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1233  (.A(\heichips25_can_lehmann_fsm/_0039_ ),
    .X(\heichips25_can_lehmann_fsm/net1232 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1234  (.A(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[1] ),
    .X(\heichips25_can_lehmann_fsm/net1233 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1235  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[15] ),
    .X(\heichips25_can_lehmann_fsm/net1234 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1236  (.A(\heichips25_can_lehmann_fsm/_0009_ ),
    .X(\heichips25_can_lehmann_fsm/net1235 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1237  (.A(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[4] ),
    .X(\heichips25_can_lehmann_fsm/net1236 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1238  (.A(\heichips25_can_lehmann_fsm/_0031_ ),
    .X(\heichips25_can_lehmann_fsm/net1237 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1239  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[22] ),
    .X(\heichips25_can_lehmann_fsm/net1238 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1240  (.A(\heichips25_can_lehmann_fsm/_0016_ ),
    .X(\heichips25_can_lehmann_fsm/net1239 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1241  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[18] ),
    .X(\heichips25_can_lehmann_fsm/net1240 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1242  (.A(\heichips25_can_lehmann_fsm/_0012_ ),
    .X(\heichips25_can_lehmann_fsm/net1241 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1243  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[9] ),
    .X(\heichips25_can_lehmann_fsm/net1242 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1244  (.A(\heichips25_can_lehmann_fsm/_0011_ ),
    .X(\heichips25_can_lehmann_fsm/net1243 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1245  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[21] ),
    .X(\heichips25_can_lehmann_fsm/net1244 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1246  (.A(\heichips25_can_lehmann_fsm/_0015_ ),
    .X(\heichips25_can_lehmann_fsm/net1245 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1247  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[20] ),
    .X(\heichips25_can_lehmann_fsm/net1246 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1248  (.A(\heichips25_can_lehmann_fsm/_0014_ ),
    .X(\heichips25_can_lehmann_fsm/net1247 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1249  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[14] ),
    .X(\heichips25_can_lehmann_fsm/net1248 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1250  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[11] ),
    .X(\heichips25_can_lehmann_fsm/net1249 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1251  (.A(\heichips25_can_lehmann_fsm/_0005_ ),
    .X(\heichips25_can_lehmann_fsm/net1250 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1252  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[16] ),
    .X(\heichips25_can_lehmann_fsm/net1251 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1253  (.A(\heichips25_can_lehmann_fsm/_0010_ ),
    .X(\heichips25_can_lehmann_fsm/net1252 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1254  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[10] ),
    .X(\heichips25_can_lehmann_fsm/net1253 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1255  (.A(\heichips25_can_lehmann_fsm/_0004_ ),
    .X(\heichips25_can_lehmann_fsm/net1254 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1256  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[0] ),
    .X(\heichips25_can_lehmann_fsm/net1255 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1257  (.A(\heichips25_can_lehmann_fsm/_0018_ ),
    .X(\heichips25_can_lehmann_fsm/net1256 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1258  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[13] ),
    .X(\heichips25_can_lehmann_fsm/net1257 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1259  (.A(\heichips25_can_lehmann_fsm/_0007_ ),
    .X(\heichips25_can_lehmann_fsm/net1258 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1260  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[19] ),
    .X(\heichips25_can_lehmann_fsm/net1259 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1261  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[12] ),
    .X(\heichips25_can_lehmann_fsm/net1260 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1262  (.A(\heichips25_can_lehmann_fsm/_0006_ ),
    .X(\heichips25_can_lehmann_fsm/net1261 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1263  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[8] ),
    .X(\heichips25_can_lehmann_fsm/net1262 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1264  (.A(\heichips25_can_lehmann_fsm/_0003_ ),
    .X(\heichips25_can_lehmann_fsm/net1263 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1265  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[4] ),
    .X(\heichips25_can_lehmann_fsm/net1264 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1266  (.A(\heichips25_can_lehmann_fsm/_0024_ ),
    .X(\heichips25_can_lehmann_fsm/net1265 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1267  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[3] ),
    .X(\heichips25_can_lehmann_fsm/net1266 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1268  (.A(\heichips25_can_lehmann_fsm/_0023_ ),
    .X(\heichips25_can_lehmann_fsm/net1267 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1269  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[7] ),
    .X(\heichips25_can_lehmann_fsm/net1268 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1270  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[1] ),
    .X(\heichips25_can_lehmann_fsm/net1269 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1271  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[5] ),
    .X(\heichips25_can_lehmann_fsm/net1270 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1272  (.A(\heichips25_can_lehmann_fsm/_0025_ ),
    .X(\heichips25_can_lehmann_fsm/net1271 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1273  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.mem_data[34] ),
    .X(\heichips25_can_lehmann_fsm/net1272 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1274  (.A(\heichips25_can_lehmann_fsm/controller.inst_mem.addr[1] ),
    .X(\heichips25_can_lehmann_fsm/net1273 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1275  (.A(\heichips25_can_lehmann_fsm/controller.alu_buffer.buffer[0] ),
    .X(\heichips25_can_lehmann_fsm/net1274 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold1276  (.A(\heichips25_sap3/sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos[0] ),
    .X(\heichips25_sap3/net1275 ));
 sg13g2_dlygate4sd3_1 \heichips25_sap3/hold1277  (.A(\heichips25_sap3/_0007_ ),
    .X(\heichips25_sap3/net1276 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1278  (.A(\heichips25_can_lehmann_fsm/controller.output_controller.keep[1] ),
    .X(\heichips25_can_lehmann_fsm/net1277 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1279  (.A(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[8] ),
    .X(\heichips25_can_lehmann_fsm/net1278 ));
 sg13g2_dlygate4sd3_1 \heichips25_can_lehmann_fsm/hold1280  (.A(\heichips25_can_lehmann_fsm/controller.counter2.counter_0[12] ),
    .X(\heichips25_can_lehmann_fsm/net1279 ));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_fill_2 FILLER_0_14 ();
 sg13g2_fill_1 FILLER_0_16 ();
 sg13g2_decap_8 FILLER_0_22 ();
 sg13g2_decap_8 FILLER_0_29 ();
 sg13g2_decap_8 FILLER_0_36 ();
 sg13g2_decap_4 FILLER_0_43 ();
 sg13g2_fill_1 FILLER_0_47 ();
 sg13g2_decap_8 FILLER_0_58 ();
 sg13g2_decap_8 FILLER_0_65 ();
 sg13g2_decap_8 FILLER_0_72 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_4 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_121 ();
 sg13g2_decap_8 FILLER_0_128 ();
 sg13g2_decap_8 FILLER_0_135 ();
 sg13g2_decap_4 FILLER_0_142 ();
 sg13g2_fill_1 FILLER_0_146 ();
 sg13g2_fill_2 FILLER_0_159 ();
 sg13g2_fill_1 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_167 ();
 sg13g2_decap_4 FILLER_0_174 ();
 sg13g2_fill_2 FILLER_0_178 ();
 sg13g2_decap_8 FILLER_0_192 ();
 sg13g2_decap_8 FILLER_0_199 ();
 sg13g2_decap_8 FILLER_0_206 ();
 sg13g2_decap_8 FILLER_0_213 ();
 sg13g2_decap_8 FILLER_0_220 ();
 sg13g2_fill_2 FILLER_0_227 ();
 sg13g2_fill_1 FILLER_0_229 ();
 sg13g2_decap_8 FILLER_0_239 ();
 sg13g2_decap_8 FILLER_0_246 ();
 sg13g2_decap_8 FILLER_0_253 ();
 sg13g2_decap_8 FILLER_0_260 ();
 sg13g2_fill_1 FILLER_0_267 ();
 sg13g2_fill_2 FILLER_0_283 ();
 sg13g2_fill_1 FILLER_0_285 ();
 sg13g2_decap_8 FILLER_0_290 ();
 sg13g2_decap_8 FILLER_0_297 ();
 sg13g2_decap_8 FILLER_0_304 ();
 sg13g2_fill_1 FILLER_0_311 ();
 sg13g2_decap_8 FILLER_0_325 ();
 sg13g2_decap_8 FILLER_0_332 ();
 sg13g2_decap_8 FILLER_0_339 ();
 sg13g2_decap_8 FILLER_0_346 ();
 sg13g2_decap_8 FILLER_0_353 ();
 sg13g2_decap_8 FILLER_0_360 ();
 sg13g2_decap_4 FILLER_0_367 ();
 sg13g2_fill_2 FILLER_0_371 ();
 sg13g2_fill_1 FILLER_0_417 ();
 sg13g2_decap_4 FILLER_0_459 ();
 sg13g2_fill_1 FILLER_0_463 ();
 sg13g2_decap_8 FILLER_0_473 ();
 sg13g2_decap_4 FILLER_0_480 ();
 sg13g2_fill_2 FILLER_0_484 ();
 sg13g2_decap_8 FILLER_0_491 ();
 sg13g2_decap_8 FILLER_0_498 ();
 sg13g2_decap_8 FILLER_0_505 ();
 sg13g2_fill_1 FILLER_0_512 ();
 sg13g2_fill_1 FILLER_0_522 ();
 sg13g2_decap_8 FILLER_0_527 ();
 sg13g2_decap_4 FILLER_0_600 ();
 sg13g2_fill_2 FILLER_0_604 ();
 sg13g2_fill_1 FILLER_0_625 ();
 sg13g2_fill_2 FILLER_0_631 ();
 sg13g2_fill_2 FILLER_0_670 ();
 sg13g2_fill_1 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_4 FILLER_0_707 ();
 sg13g2_fill_2 FILLER_0_711 ();
 sg13g2_fill_1 FILLER_0_745 ();
 sg13g2_decap_4 FILLER_0_755 ();
 sg13g2_fill_1 FILLER_0_759 ();
 sg13g2_decap_4 FILLER_0_787 ();
 sg13g2_fill_1 FILLER_0_791 ();
 sg13g2_fill_2 FILLER_0_824 ();
 sg13g2_fill_2 FILLER_0_831 ();
 sg13g2_fill_2 FILLER_0_838 ();
 sg13g2_fill_1 FILLER_0_840 ();
 sg13g2_decap_4 FILLER_0_846 ();
 sg13g2_fill_2 FILLER_0_850 ();
 sg13g2_fill_1 FILLER_0_873 ();
 sg13g2_decap_8 FILLER_0_901 ();
 sg13g2_decap_8 FILLER_0_908 ();
 sg13g2_decap_8 FILLER_0_915 ();
 sg13g2_decap_8 FILLER_0_922 ();
 sg13g2_decap_8 FILLER_0_929 ();
 sg13g2_decap_8 FILLER_0_936 ();
 sg13g2_decap_8 FILLER_0_943 ();
 sg13g2_decap_8 FILLER_0_950 ();
 sg13g2_decap_8 FILLER_0_957 ();
 sg13g2_decap_8 FILLER_0_964 ();
 sg13g2_decap_8 FILLER_0_971 ();
 sg13g2_decap_8 FILLER_0_978 ();
 sg13g2_decap_8 FILLER_0_985 ();
 sg13g2_decap_8 FILLER_0_992 ();
 sg13g2_decap_8 FILLER_0_999 ();
 sg13g2_decap_8 FILLER_0_1006 ();
 sg13g2_decap_8 FILLER_0_1013 ();
 sg13g2_decap_8 FILLER_0_1020 ();
 sg13g2_fill_2 FILLER_0_1027 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_fill_2 FILLER_1_7 ();
 sg13g2_decap_4 FILLER_1_33 ();
 sg13g2_decap_8 FILLER_1_68 ();
 sg13g2_decap_4 FILLER_1_93 ();
 sg13g2_fill_1 FILLER_1_97 ();
 sg13g2_fill_2 FILLER_1_117 ();
 sg13g2_fill_1 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_125 ();
 sg13g2_decap_8 FILLER_1_132 ();
 sg13g2_fill_1 FILLER_1_139 ();
 sg13g2_fill_1 FILLER_1_153 ();
 sg13g2_fill_2 FILLER_1_174 ();
 sg13g2_decap_8 FILLER_1_205 ();
 sg13g2_fill_2 FILLER_1_212 ();
 sg13g2_fill_1 FILLER_1_214 ();
 sg13g2_fill_2 FILLER_1_267 ();
 sg13g2_fill_1 FILLER_1_269 ();
 sg13g2_fill_2 FILLER_1_276 ();
 sg13g2_fill_1 FILLER_1_278 ();
 sg13g2_fill_2 FILLER_1_316 ();
 sg13g2_fill_1 FILLER_1_345 ();
 sg13g2_fill_2 FILLER_1_511 ();
 sg13g2_decap_4 FILLER_1_540 ();
 sg13g2_decap_4 FILLER_1_571 ();
 sg13g2_fill_1 FILLER_1_636 ();
 sg13g2_fill_2 FILLER_1_669 ();
 sg13g2_fill_1 FILLER_1_671 ();
 sg13g2_fill_2 FILLER_1_699 ();
 sg13g2_fill_1 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_912 ();
 sg13g2_decap_8 FILLER_1_919 ();
 sg13g2_decap_8 FILLER_1_926 ();
 sg13g2_decap_8 FILLER_1_933 ();
 sg13g2_decap_8 FILLER_1_940 ();
 sg13g2_decap_8 FILLER_1_947 ();
 sg13g2_decap_8 FILLER_1_954 ();
 sg13g2_decap_8 FILLER_1_961 ();
 sg13g2_decap_8 FILLER_1_968 ();
 sg13g2_decap_8 FILLER_1_975 ();
 sg13g2_decap_8 FILLER_1_982 ();
 sg13g2_decap_8 FILLER_1_989 ();
 sg13g2_decap_8 FILLER_1_996 ();
 sg13g2_decap_8 FILLER_1_1003 ();
 sg13g2_decap_8 FILLER_1_1010 ();
 sg13g2_decap_8 FILLER_1_1017 ();
 sg13g2_decap_4 FILLER_1_1024 ();
 sg13g2_fill_1 FILLER_1_1028 ();
 sg13g2_decap_8 FILLER_2_4 ();
 sg13g2_decap_4 FILLER_2_11 ();
 sg13g2_fill_1 FILLER_2_15 ();
 sg13g2_fill_2 FILLER_2_30 ();
 sg13g2_decap_8 FILLER_2_60 ();
 sg13g2_decap_8 FILLER_2_67 ();
 sg13g2_decap_4 FILLER_2_74 ();
 sg13g2_fill_1 FILLER_2_78 ();
 sg13g2_fill_1 FILLER_2_89 ();
 sg13g2_fill_2 FILLER_2_109 ();
 sg13g2_fill_1 FILLER_2_111 ();
 sg13g2_decap_8 FILLER_2_117 ();
 sg13g2_fill_1 FILLER_2_124 ();
 sg13g2_decap_8 FILLER_2_135 ();
 sg13g2_decap_4 FILLER_2_158 ();
 sg13g2_fill_1 FILLER_2_162 ();
 sg13g2_fill_2 FILLER_2_168 ();
 sg13g2_fill_1 FILLER_2_170 ();
 sg13g2_fill_2 FILLER_2_180 ();
 sg13g2_fill_1 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_193 ();
 sg13g2_decap_8 FILLER_2_200 ();
 sg13g2_fill_1 FILLER_2_207 ();
 sg13g2_fill_2 FILLER_2_219 ();
 sg13g2_fill_1 FILLER_2_221 ();
 sg13g2_fill_1 FILLER_2_226 ();
 sg13g2_decap_8 FILLER_2_239 ();
 sg13g2_decap_8 FILLER_2_246 ();
 sg13g2_decap_8 FILLER_2_253 ();
 sg13g2_fill_1 FILLER_2_260 ();
 sg13g2_decap_8 FILLER_2_284 ();
 sg13g2_fill_1 FILLER_2_291 ();
 sg13g2_fill_1 FILLER_2_324 ();
 sg13g2_decap_8 FILLER_2_333 ();
 sg13g2_decap_8 FILLER_2_340 ();
 sg13g2_decap_4 FILLER_2_347 ();
 sg13g2_decap_8 FILLER_2_382 ();
 sg13g2_decap_8 FILLER_2_389 ();
 sg13g2_decap_8 FILLER_2_396 ();
 sg13g2_decap_8 FILLER_2_403 ();
 sg13g2_fill_2 FILLER_2_410 ();
 sg13g2_decap_8 FILLER_2_416 ();
 sg13g2_fill_2 FILLER_2_423 ();
 sg13g2_fill_1 FILLER_2_425 ();
 sg13g2_decap_8 FILLER_2_436 ();
 sg13g2_decap_8 FILLER_2_443 ();
 sg13g2_decap_8 FILLER_2_450 ();
 sg13g2_decap_4 FILLER_2_457 ();
 sg13g2_fill_2 FILLER_2_461 ();
 sg13g2_decap_4 FILLER_2_475 ();
 sg13g2_fill_2 FILLER_2_479 ();
 sg13g2_decap_4 FILLER_2_490 ();
 sg13g2_fill_1 FILLER_2_494 ();
 sg13g2_decap_8 FILLER_2_507 ();
 sg13g2_fill_1 FILLER_2_514 ();
 sg13g2_decap_8 FILLER_2_519 ();
 sg13g2_fill_2 FILLER_2_526 ();
 sg13g2_decap_4 FILLER_2_606 ();
 sg13g2_fill_1 FILLER_2_643 ();
 sg13g2_fill_1 FILLER_2_663 ();
 sg13g2_decap_8 FILLER_2_730 ();
 sg13g2_fill_2 FILLER_2_737 ();
 sg13g2_decap_4 FILLER_2_744 ();
 sg13g2_fill_2 FILLER_2_753 ();
 sg13g2_fill_1 FILLER_2_755 ();
 sg13g2_decap_8 FILLER_2_765 ();
 sg13g2_decap_8 FILLER_2_772 ();
 sg13g2_decap_8 FILLER_2_784 ();
 sg13g2_fill_2 FILLER_2_791 ();
 sg13g2_fill_1 FILLER_2_797 ();
 sg13g2_fill_2 FILLER_2_810 ();
 sg13g2_fill_2 FILLER_2_842 ();
 sg13g2_decap_4 FILLER_2_853 ();
 sg13g2_fill_1 FILLER_2_857 ();
 sg13g2_fill_2 FILLER_2_868 ();
 sg13g2_fill_2 FILLER_2_884 ();
 sg13g2_fill_1 FILLER_2_903 ();
 sg13g2_decap_8 FILLER_2_913 ();
 sg13g2_decap_8 FILLER_2_920 ();
 sg13g2_decap_8 FILLER_2_930 ();
 sg13g2_decap_8 FILLER_2_937 ();
 sg13g2_decap_8 FILLER_2_944 ();
 sg13g2_decap_8 FILLER_2_951 ();
 sg13g2_decap_8 FILLER_2_958 ();
 sg13g2_decap_8 FILLER_2_965 ();
 sg13g2_decap_8 FILLER_2_972 ();
 sg13g2_decap_8 FILLER_2_979 ();
 sg13g2_decap_8 FILLER_2_986 ();
 sg13g2_decap_8 FILLER_2_993 ();
 sg13g2_decap_8 FILLER_2_1000 ();
 sg13g2_decap_8 FILLER_2_1007 ();
 sg13g2_decap_8 FILLER_2_1014 ();
 sg13g2_decap_8 FILLER_2_1021 ();
 sg13g2_fill_1 FILLER_2_1028 ();
 sg13g2_decap_8 FILLER_3_4 ();
 sg13g2_decap_4 FILLER_3_11 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_58 ();
 sg13g2_fill_1 FILLER_3_65 ();
 sg13g2_decap_4 FILLER_3_77 ();
 sg13g2_fill_2 FILLER_3_81 ();
 sg13g2_decap_8 FILLER_3_88 ();
 sg13g2_decap_8 FILLER_3_95 ();
 sg13g2_decap_4 FILLER_3_102 ();
 sg13g2_decap_8 FILLER_3_111 ();
 sg13g2_decap_4 FILLER_3_118 ();
 sg13g2_fill_2 FILLER_3_132 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_fill_2 FILLER_3_168 ();
 sg13g2_fill_1 FILLER_3_170 ();
 sg13g2_decap_4 FILLER_3_175 ();
 sg13g2_fill_1 FILLER_3_179 ();
 sg13g2_fill_2 FILLER_3_188 ();
 sg13g2_decap_8 FILLER_3_195 ();
 sg13g2_fill_2 FILLER_3_202 ();
 sg13g2_decap_8 FILLER_3_209 ();
 sg13g2_fill_2 FILLER_3_216 ();
 sg13g2_fill_2 FILLER_3_231 ();
 sg13g2_fill_1 FILLER_3_233 ();
 sg13g2_fill_2 FILLER_3_243 ();
 sg13g2_fill_1 FILLER_3_245 ();
 sg13g2_fill_2 FILLER_3_254 ();
 sg13g2_fill_1 FILLER_3_256 ();
 sg13g2_fill_2 FILLER_3_269 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_fill_1 FILLER_3_294 ();
 sg13g2_decap_4 FILLER_3_319 ();
 sg13g2_decap_8 FILLER_3_327 ();
 sg13g2_decap_8 FILLER_3_334 ();
 sg13g2_fill_1 FILLER_3_341 ();
 sg13g2_decap_4 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_366 ();
 sg13g2_fill_2 FILLER_3_373 ();
 sg13g2_fill_1 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_397 ();
 sg13g2_fill_2 FILLER_3_404 ();
 sg13g2_fill_1 FILLER_3_419 ();
 sg13g2_decap_4 FILLER_3_430 ();
 sg13g2_fill_1 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_440 ();
 sg13g2_decap_8 FILLER_3_456 ();
 sg13g2_fill_2 FILLER_3_463 ();
 sg13g2_decap_8 FILLER_3_478 ();
 sg13g2_decap_8 FILLER_3_485 ();
 sg13g2_decap_8 FILLER_3_492 ();
 sg13g2_fill_2 FILLER_3_499 ();
 sg13g2_fill_1 FILLER_3_501 ();
 sg13g2_decap_8 FILLER_3_518 ();
 sg13g2_fill_2 FILLER_3_525 ();
 sg13g2_decap_4 FILLER_3_544 ();
 sg13g2_decap_4 FILLER_3_557 ();
 sg13g2_decap_8 FILLER_3_574 ();
 sg13g2_decap_4 FILLER_3_585 ();
 sg13g2_fill_1 FILLER_3_589 ();
 sg13g2_decap_4 FILLER_3_621 ();
 sg13g2_fill_2 FILLER_3_625 ();
 sg13g2_decap_4 FILLER_3_631 ();
 sg13g2_fill_2 FILLER_3_662 ();
 sg13g2_fill_1 FILLER_3_664 ();
 sg13g2_decap_4 FILLER_3_696 ();
 sg13g2_decap_8 FILLER_3_722 ();
 sg13g2_fill_2 FILLER_3_729 ();
 sg13g2_fill_1 FILLER_3_731 ();
 sg13g2_fill_1 FILLER_3_764 ();
 sg13g2_decap_8 FILLER_3_783 ();
 sg13g2_fill_1 FILLER_3_790 ();
 sg13g2_fill_1 FILLER_3_800 ();
 sg13g2_decap_4 FILLER_3_804 ();
 sg13g2_decap_4 FILLER_3_850 ();
 sg13g2_fill_2 FILLER_3_854 ();
 sg13g2_fill_2 FILLER_3_883 ();
 sg13g2_fill_1 FILLER_3_885 ();
 sg13g2_fill_2 FILLER_3_913 ();
 sg13g2_fill_1 FILLER_3_924 ();
 sg13g2_fill_2 FILLER_3_944 ();
 sg13g2_fill_1 FILLER_3_946 ();
 sg13g2_decap_8 FILLER_3_956 ();
 sg13g2_decap_8 FILLER_3_963 ();
 sg13g2_decap_8 FILLER_3_970 ();
 sg13g2_decap_8 FILLER_3_977 ();
 sg13g2_decap_8 FILLER_3_984 ();
 sg13g2_decap_8 FILLER_3_991 ();
 sg13g2_decap_8 FILLER_3_998 ();
 sg13g2_decap_8 FILLER_3_1005 ();
 sg13g2_decap_8 FILLER_3_1012 ();
 sg13g2_decap_8 FILLER_3_1019 ();
 sg13g2_fill_2 FILLER_3_1026 ();
 sg13g2_fill_1 FILLER_3_1028 ();
 sg13g2_fill_1 FILLER_4_4 ();
 sg13g2_fill_1 FILLER_4_26 ();
 sg13g2_decap_4 FILLER_4_37 ();
 sg13g2_decap_8 FILLER_4_46 ();
 sg13g2_decap_8 FILLER_4_53 ();
 sg13g2_decap_8 FILLER_4_60 ();
 sg13g2_fill_1 FILLER_4_67 ();
 sg13g2_fill_1 FILLER_4_79 ();
 sg13g2_decap_8 FILLER_4_92 ();
 sg13g2_decap_4 FILLER_4_99 ();
 sg13g2_fill_2 FILLER_4_103 ();
 sg13g2_fill_1 FILLER_4_110 ();
 sg13g2_decap_8 FILLER_4_116 ();
 sg13g2_decap_8 FILLER_4_123 ();
 sg13g2_decap_8 FILLER_4_130 ();
 sg13g2_fill_2 FILLER_4_137 ();
 sg13g2_fill_2 FILLER_4_147 ();
 sg13g2_fill_1 FILLER_4_149 ();
 sg13g2_decap_8 FILLER_4_160 ();
 sg13g2_fill_2 FILLER_4_167 ();
 sg13g2_decap_4 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_fill_2 FILLER_4_210 ();
 sg13g2_fill_2 FILLER_4_221 ();
 sg13g2_decap_8 FILLER_4_227 ();
 sg13g2_fill_1 FILLER_4_234 ();
 sg13g2_decap_4 FILLER_4_255 ();
 sg13g2_decap_8 FILLER_4_264 ();
 sg13g2_fill_2 FILLER_4_271 ();
 sg13g2_fill_1 FILLER_4_285 ();
 sg13g2_decap_4 FILLER_4_290 ();
 sg13g2_decap_8 FILLER_4_299 ();
 sg13g2_decap_4 FILLER_4_306 ();
 sg13g2_fill_2 FILLER_4_310 ();
 sg13g2_fill_1 FILLER_4_317 ();
 sg13g2_fill_1 FILLER_4_323 ();
 sg13g2_fill_2 FILLER_4_338 ();
 sg13g2_fill_1 FILLER_4_352 ();
 sg13g2_decap_4 FILLER_4_358 ();
 sg13g2_fill_1 FILLER_4_362 ();
 sg13g2_fill_2 FILLER_4_385 ();
 sg13g2_fill_1 FILLER_4_387 ();
 sg13g2_fill_2 FILLER_4_393 ();
 sg13g2_fill_2 FILLER_4_438 ();
 sg13g2_fill_2 FILLER_4_452 ();
 sg13g2_decap_4 FILLER_4_459 ();
 sg13g2_fill_2 FILLER_4_478 ();
 sg13g2_fill_2 FILLER_4_492 ();
 sg13g2_fill_1 FILLER_4_506 ();
 sg13g2_fill_2 FILLER_4_523 ();
 sg13g2_fill_1 FILLER_4_525 ();
 sg13g2_decap_8 FILLER_4_544 ();
 sg13g2_fill_2 FILLER_4_551 ();
 sg13g2_fill_1 FILLER_4_553 ();
 sg13g2_fill_1 FILLER_4_606 ();
 sg13g2_fill_2 FILLER_4_625 ();
 sg13g2_fill_1 FILLER_4_645 ();
 sg13g2_fill_2 FILLER_4_655 ();
 sg13g2_fill_2 FILLER_4_675 ();
 sg13g2_fill_1 FILLER_4_690 ();
 sg13g2_fill_1 FILLER_4_737 ();
 sg13g2_fill_2 FILLER_4_760 ();
 sg13g2_decap_4 FILLER_4_831 ();
 sg13g2_decap_8 FILLER_4_847 ();
 sg13g2_decap_8 FILLER_4_854 ();
 sg13g2_decap_8 FILLER_4_870 ();
 sg13g2_decap_8 FILLER_4_877 ();
 sg13g2_fill_1 FILLER_4_884 ();
 sg13g2_fill_1 FILLER_4_890 ();
 sg13g2_fill_2 FILLER_4_895 ();
 sg13g2_fill_1 FILLER_4_959 ();
 sg13g2_fill_2 FILLER_4_964 ();
 sg13g2_decap_8 FILLER_4_980 ();
 sg13g2_decap_8 FILLER_4_987 ();
 sg13g2_decap_8 FILLER_4_994 ();
 sg13g2_decap_8 FILLER_4_1001 ();
 sg13g2_decap_8 FILLER_4_1008 ();
 sg13g2_decap_8 FILLER_4_1015 ();
 sg13g2_decap_8 FILLER_4_1022 ();
 sg13g2_decap_8 FILLER_5_4 ();
 sg13g2_fill_1 FILLER_5_11 ();
 sg13g2_fill_1 FILLER_5_37 ();
 sg13g2_fill_1 FILLER_5_43 ();
 sg13g2_decap_8 FILLER_5_66 ();
 sg13g2_fill_1 FILLER_5_73 ();
 sg13g2_fill_2 FILLER_5_78 ();
 sg13g2_decap_4 FILLER_5_91 ();
 sg13g2_fill_1 FILLER_5_95 ();
 sg13g2_decap_4 FILLER_5_102 ();
 sg13g2_fill_1 FILLER_5_109 ();
 sg13g2_fill_1 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_129 ();
 sg13g2_decap_8 FILLER_5_136 ();
 sg13g2_fill_2 FILLER_5_143 ();
 sg13g2_fill_1 FILLER_5_145 ();
 sg13g2_decap_8 FILLER_5_162 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_fill_2 FILLER_5_203 ();
 sg13g2_fill_1 FILLER_5_221 ();
 sg13g2_fill_1 FILLER_5_226 ();
 sg13g2_fill_2 FILLER_5_231 ();
 sg13g2_fill_1 FILLER_5_233 ();
 sg13g2_decap_8 FILLER_5_240 ();
 sg13g2_decap_8 FILLER_5_247 ();
 sg13g2_decap_4 FILLER_5_254 ();
 sg13g2_fill_1 FILLER_5_258 ();
 sg13g2_decap_8 FILLER_5_267 ();
 sg13g2_decap_4 FILLER_5_274 ();
 sg13g2_fill_2 FILLER_5_292 ();
 sg13g2_fill_1 FILLER_5_294 ();
 sg13g2_fill_2 FILLER_5_315 ();
 sg13g2_decap_4 FILLER_5_325 ();
 sg13g2_fill_2 FILLER_5_351 ();
 sg13g2_fill_1 FILLER_5_353 ();
 sg13g2_decap_8 FILLER_5_394 ();
 sg13g2_fill_2 FILLER_5_401 ();
 sg13g2_decap_4 FILLER_5_421 ();
 sg13g2_fill_2 FILLER_5_425 ();
 sg13g2_decap_8 FILLER_5_448 ();
 sg13g2_decap_8 FILLER_5_455 ();
 sg13g2_decap_4 FILLER_5_462 ();
 sg13g2_fill_2 FILLER_5_466 ();
 sg13g2_decap_4 FILLER_5_486 ();
 sg13g2_fill_1 FILLER_5_490 ();
 sg13g2_decap_4 FILLER_5_509 ();
 sg13g2_fill_2 FILLER_5_523 ();
 sg13g2_decap_4 FILLER_5_554 ();
 sg13g2_fill_2 FILLER_5_558 ();
 sg13g2_fill_1 FILLER_5_577 ();
 sg13g2_fill_1 FILLER_5_610 ();
 sg13g2_fill_2 FILLER_5_714 ();
 sg13g2_fill_1 FILLER_5_716 ();
 sg13g2_fill_2 FILLER_5_728 ();
 sg13g2_fill_1 FILLER_5_730 ();
 sg13g2_decap_8 FILLER_5_769 ();
 sg13g2_decap_8 FILLER_5_781 ();
 sg13g2_fill_2 FILLER_5_788 ();
 sg13g2_fill_2 FILLER_5_799 ();
 sg13g2_fill_2 FILLER_5_804 ();
 sg13g2_fill_1 FILLER_5_806 ();
 sg13g2_decap_8 FILLER_5_833 ();
 sg13g2_fill_2 FILLER_5_840 ();
 sg13g2_fill_1 FILLER_5_842 ();
 sg13g2_fill_2 FILLER_5_861 ();
 sg13g2_fill_1 FILLER_5_863 ();
 sg13g2_fill_2 FILLER_5_869 ();
 sg13g2_decap_8 FILLER_5_877 ();
 sg13g2_fill_2 FILLER_5_887 ();
 sg13g2_decap_4 FILLER_5_901 ();
 sg13g2_fill_2 FILLER_5_924 ();
 sg13g2_fill_1 FILLER_5_932 ();
 sg13g2_fill_2 FILLER_5_938 ();
 sg13g2_fill_2 FILLER_5_967 ();
 sg13g2_decap_8 FILLER_5_996 ();
 sg13g2_decap_8 FILLER_5_1003 ();
 sg13g2_decap_8 FILLER_5_1010 ();
 sg13g2_decap_8 FILLER_5_1017 ();
 sg13g2_decap_4 FILLER_5_1024 ();
 sg13g2_fill_1 FILLER_5_1028 ();
 sg13g2_decap_8 FILLER_6_4 ();
 sg13g2_decap_8 FILLER_6_34 ();
 sg13g2_decap_8 FILLER_6_41 ();
 sg13g2_decap_8 FILLER_6_48 ();
 sg13g2_decap_4 FILLER_6_55 ();
 sg13g2_fill_1 FILLER_6_59 ();
 sg13g2_fill_2 FILLER_6_65 ();
 sg13g2_fill_1 FILLER_6_67 ();
 sg13g2_decap_8 FILLER_6_72 ();
 sg13g2_fill_2 FILLER_6_83 ();
 sg13g2_decap_4 FILLER_6_89 ();
 sg13g2_decap_8 FILLER_6_97 ();
 sg13g2_decap_8 FILLER_6_104 ();
 sg13g2_fill_2 FILLER_6_111 ();
 sg13g2_decap_4 FILLER_6_122 ();
 sg13g2_decap_8 FILLER_6_132 ();
 sg13g2_decap_8 FILLER_6_139 ();
 sg13g2_decap_4 FILLER_6_146 ();
 sg13g2_decap_8 FILLER_6_160 ();
 sg13g2_fill_2 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_183 ();
 sg13g2_decap_4 FILLER_6_190 ();
 sg13g2_fill_2 FILLER_6_194 ();
 sg13g2_decap_8 FILLER_6_207 ();
 sg13g2_fill_2 FILLER_6_214 ();
 sg13g2_fill_1 FILLER_6_216 ();
 sg13g2_decap_8 FILLER_6_225 ();
 sg13g2_decap_4 FILLER_6_247 ();
 sg13g2_fill_2 FILLER_6_255 ();
 sg13g2_decap_8 FILLER_6_274 ();
 sg13g2_decap_8 FILLER_6_281 ();
 sg13g2_decap_4 FILLER_6_288 ();
 sg13g2_fill_2 FILLER_6_292 ();
 sg13g2_decap_4 FILLER_6_298 ();
 sg13g2_fill_1 FILLER_6_302 ();
 sg13g2_decap_8 FILLER_6_310 ();
 sg13g2_decap_8 FILLER_6_317 ();
 sg13g2_decap_8 FILLER_6_324 ();
 sg13g2_fill_2 FILLER_6_331 ();
 sg13g2_fill_1 FILLER_6_338 ();
 sg13g2_fill_2 FILLER_6_360 ();
 sg13g2_fill_2 FILLER_6_366 ();
 sg13g2_fill_1 FILLER_6_368 ();
 sg13g2_fill_2 FILLER_6_377 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_4 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_405 ();
 sg13g2_decap_8 FILLER_6_412 ();
 sg13g2_decap_8 FILLER_6_419 ();
 sg13g2_decap_8 FILLER_6_426 ();
 sg13g2_decap_4 FILLER_6_433 ();
 sg13g2_fill_1 FILLER_6_437 ();
 sg13g2_fill_2 FILLER_6_443 ();
 sg13g2_fill_1 FILLER_6_445 ();
 sg13g2_decap_8 FILLER_6_456 ();
 sg13g2_decap_8 FILLER_6_463 ();
 sg13g2_decap_8 FILLER_6_470 ();
 sg13g2_fill_2 FILLER_6_477 ();
 sg13g2_fill_1 FILLER_6_479 ();
 sg13g2_decap_8 FILLER_6_489 ();
 sg13g2_decap_4 FILLER_6_496 ();
 sg13g2_fill_2 FILLER_6_500 ();
 sg13g2_decap_8 FILLER_6_510 ();
 sg13g2_decap_8 FILLER_6_517 ();
 sg13g2_decap_8 FILLER_6_524 ();
 sg13g2_fill_2 FILLER_6_531 ();
 sg13g2_fill_2 FILLER_6_543 ();
 sg13g2_fill_1 FILLER_6_545 ();
 sg13g2_decap_4 FILLER_6_551 ();
 sg13g2_decap_4 FILLER_6_560 ();
 sg13g2_fill_2 FILLER_6_593 ();
 sg13g2_fill_1 FILLER_6_595 ();
 sg13g2_decap_4 FILLER_6_633 ();
 sg13g2_fill_2 FILLER_6_637 ();
 sg13g2_fill_2 FILLER_6_674 ();
 sg13g2_fill_1 FILLER_6_693 ();
 sg13g2_fill_2 FILLER_6_725 ();
 sg13g2_fill_1 FILLER_6_727 ();
 sg13g2_fill_1 FILLER_6_758 ();
 sg13g2_decap_8 FILLER_6_778 ();
 sg13g2_fill_1 FILLER_6_785 ();
 sg13g2_fill_1 FILLER_6_826 ();
 sg13g2_fill_2 FILLER_6_838 ();
 sg13g2_fill_1 FILLER_6_867 ();
 sg13g2_fill_1 FILLER_6_963 ();
 sg13g2_decap_4 FILLER_6_996 ();
 sg13g2_fill_1 FILLER_6_1000 ();
 sg13g2_fill_2 FILLER_6_1006 ();
 sg13g2_fill_2 FILLER_6_1012 ();
 sg13g2_fill_1 FILLER_6_1014 ();
 sg13g2_decap_4 FILLER_6_1024 ();
 sg13g2_fill_1 FILLER_6_1028 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_fill_2 FILLER_7_7 ();
 sg13g2_fill_1 FILLER_7_9 ();
 sg13g2_fill_2 FILLER_7_42 ();
 sg13g2_fill_1 FILLER_7_44 ();
 sg13g2_decap_8 FILLER_7_51 ();
 sg13g2_decap_8 FILLER_7_58 ();
 sg13g2_decap_4 FILLER_7_65 ();
 sg13g2_fill_1 FILLER_7_69 ();
 sg13g2_decap_8 FILLER_7_79 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_4 FILLER_7_98 ();
 sg13g2_fill_2 FILLER_7_102 ();
 sg13g2_fill_2 FILLER_7_109 ();
 sg13g2_fill_2 FILLER_7_116 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_4 FILLER_7_140 ();
 sg13g2_fill_1 FILLER_7_144 ();
 sg13g2_fill_1 FILLER_7_149 ();
 sg13g2_fill_2 FILLER_7_155 ();
 sg13g2_decap_4 FILLER_7_166 ();
 sg13g2_fill_2 FILLER_7_170 ();
 sg13g2_decap_4 FILLER_7_184 ();
 sg13g2_fill_1 FILLER_7_188 ();
 sg13g2_decap_8 FILLER_7_207 ();
 sg13g2_decap_8 FILLER_7_214 ();
 sg13g2_decap_8 FILLER_7_226 ();
 sg13g2_fill_1 FILLER_7_233 ();
 sg13g2_decap_8 FILLER_7_243 ();
 sg13g2_decap_8 FILLER_7_250 ();
 sg13g2_decap_4 FILLER_7_257 ();
 sg13g2_fill_1 FILLER_7_261 ();
 sg13g2_decap_8 FILLER_7_276 ();
 sg13g2_fill_2 FILLER_7_283 ();
 sg13g2_fill_1 FILLER_7_285 ();
 sg13g2_decap_4 FILLER_7_290 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_4 FILLER_7_329 ();
 sg13g2_fill_2 FILLER_7_333 ();
 sg13g2_decap_8 FILLER_7_349 ();
 sg13g2_decap_8 FILLER_7_356 ();
 sg13g2_decap_8 FILLER_7_363 ();
 sg13g2_decap_4 FILLER_7_370 ();
 sg13g2_fill_2 FILLER_7_386 ();
 sg13g2_decap_4 FILLER_7_404 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_4 FILLER_7_416 ();
 sg13g2_fill_2 FILLER_7_430 ();
 sg13g2_fill_1 FILLER_7_432 ();
 sg13g2_decap_4 FILLER_7_443 ();
 sg13g2_fill_2 FILLER_7_447 ();
 sg13g2_decap_4 FILLER_7_458 ();
 sg13g2_fill_1 FILLER_7_462 ();
 sg13g2_decap_8 FILLER_7_469 ();
 sg13g2_decap_8 FILLER_7_488 ();
 sg13g2_decap_4 FILLER_7_495 ();
 sg13g2_fill_2 FILLER_7_499 ();
 sg13g2_fill_2 FILLER_7_511 ();
 sg13g2_decap_8 FILLER_7_521 ();
 sg13g2_decap_8 FILLER_7_528 ();
 sg13g2_fill_1 FILLER_7_535 ();
 sg13g2_fill_1 FILLER_7_550 ();
 sg13g2_fill_2 FILLER_7_586 ();
 sg13g2_fill_1 FILLER_7_624 ();
 sg13g2_fill_2 FILLER_7_715 ();
 sg13g2_fill_2 FILLER_7_731 ();
 sg13g2_decap_4 FILLER_7_743 ();
 sg13g2_fill_2 FILLER_7_761 ();
 sg13g2_decap_8 FILLER_7_784 ();
 sg13g2_decap_8 FILLER_7_795 ();
 sg13g2_fill_1 FILLER_7_802 ();
 sg13g2_fill_2 FILLER_7_823 ();
 sg13g2_fill_1 FILLER_7_825 ();
 sg13g2_decap_4 FILLER_7_837 ();
 sg13g2_fill_2 FILLER_7_841 ();
 sg13g2_fill_2 FILLER_7_852 ();
 sg13g2_fill_1 FILLER_7_854 ();
 sg13g2_decap_8 FILLER_7_888 ();
 sg13g2_fill_1 FILLER_7_895 ();
 sg13g2_decap_8 FILLER_7_899 ();
 sg13g2_decap_4 FILLER_7_938 ();
 sg13g2_fill_1 FILLER_7_969 ();
 sg13g2_fill_2 FILLER_7_1000 ();
 sg13g2_decap_8 FILLER_8_4 ();
 sg13g2_decap_4 FILLER_8_11 ();
 sg13g2_decap_8 FILLER_8_25 ();
 sg13g2_decap_8 FILLER_8_32 ();
 sg13g2_decap_8 FILLER_8_39 ();
 sg13g2_fill_2 FILLER_8_46 ();
 sg13g2_decap_8 FILLER_8_65 ();
 sg13g2_decap_8 FILLER_8_72 ();
 sg13g2_fill_2 FILLER_8_88 ();
 sg13g2_decap_8 FILLER_8_99 ();
 sg13g2_decap_4 FILLER_8_106 ();
 sg13g2_fill_1 FILLER_8_110 ();
 sg13g2_decap_4 FILLER_8_117 ();
 sg13g2_fill_1 FILLER_8_121 ();
 sg13g2_fill_2 FILLER_8_126 ();
 sg13g2_fill_1 FILLER_8_128 ();
 sg13g2_fill_2 FILLER_8_139 ();
 sg13g2_fill_2 FILLER_8_151 ();
 sg13g2_decap_4 FILLER_8_158 ();
 sg13g2_fill_2 FILLER_8_162 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_4 FILLER_8_175 ();
 sg13g2_fill_1 FILLER_8_179 ();
 sg13g2_decap_8 FILLER_8_184 ();
 sg13g2_decap_4 FILLER_8_191 ();
 sg13g2_fill_2 FILLER_8_195 ();
 sg13g2_fill_2 FILLER_8_201 ();
 sg13g2_fill_1 FILLER_8_203 ();
 sg13g2_fill_2 FILLER_8_223 ();
 sg13g2_fill_1 FILLER_8_225 ();
 sg13g2_fill_2 FILLER_8_237 ();
 sg13g2_fill_1 FILLER_8_239 ();
 sg13g2_decap_4 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_279 ();
 sg13g2_fill_2 FILLER_8_286 ();
 sg13g2_decap_4 FILLER_8_292 ();
 sg13g2_fill_1 FILLER_8_296 ();
 sg13g2_fill_2 FILLER_8_307 ();
 sg13g2_decap_8 FILLER_8_318 ();
 sg13g2_fill_1 FILLER_8_325 ();
 sg13g2_fill_1 FILLER_8_334 ();
 sg13g2_decap_8 FILLER_8_344 ();
 sg13g2_decap_8 FILLER_8_351 ();
 sg13g2_decap_4 FILLER_8_358 ();
 sg13g2_decap_8 FILLER_8_386 ();
 sg13g2_decap_8 FILLER_8_393 ();
 sg13g2_fill_1 FILLER_8_411 ();
 sg13g2_decap_8 FILLER_8_416 ();
 sg13g2_decap_8 FILLER_8_423 ();
 sg13g2_fill_2 FILLER_8_430 ();
 sg13g2_fill_1 FILLER_8_432 ();
 sg13g2_decap_8 FILLER_8_444 ();
 sg13g2_decap_8 FILLER_8_451 ();
 sg13g2_decap_8 FILLER_8_458 ();
 sg13g2_decap_8 FILLER_8_470 ();
 sg13g2_decap_4 FILLER_8_477 ();
 sg13g2_fill_1 FILLER_8_481 ();
 sg13g2_decap_4 FILLER_8_488 ();
 sg13g2_fill_2 FILLER_8_492 ();
 sg13g2_decap_8 FILLER_8_524 ();
 sg13g2_decap_8 FILLER_8_531 ();
 sg13g2_decap_8 FILLER_8_538 ();
 sg13g2_fill_2 FILLER_8_555 ();
 sg13g2_decap_8 FILLER_8_588 ();
 sg13g2_fill_1 FILLER_8_595 ();
 sg13g2_decap_4 FILLER_8_600 ();
 sg13g2_fill_1 FILLER_8_604 ();
 sg13g2_fill_2 FILLER_8_642 ();
 sg13g2_decap_8 FILLER_8_689 ();
 sg13g2_decap_4 FILLER_8_696 ();
 sg13g2_fill_2 FILLER_8_704 ();
 sg13g2_fill_1 FILLER_8_711 ();
 sg13g2_decap_4 FILLER_8_777 ();
 sg13g2_decap_4 FILLER_8_804 ();
 sg13g2_fill_1 FILLER_8_808 ();
 sg13g2_decap_4 FILLER_8_841 ();
 sg13g2_fill_1 FILLER_8_845 ();
 sg13g2_fill_2 FILLER_8_855 ();
 sg13g2_fill_2 FILLER_8_871 ();
 sg13g2_fill_2 FILLER_8_879 ();
 sg13g2_decap_8 FILLER_8_952 ();
 sg13g2_decap_4 FILLER_8_959 ();
 sg13g2_fill_1 FILLER_8_963 ();
 sg13g2_fill_2 FILLER_8_986 ();
 sg13g2_decap_4 FILLER_8_1024 ();
 sg13g2_fill_1 FILLER_8_1028 ();
 sg13g2_decap_8 FILLER_9_8 ();
 sg13g2_fill_2 FILLER_9_15 ();
 sg13g2_fill_2 FILLER_9_26 ();
 sg13g2_decap_8 FILLER_9_38 ();
 sg13g2_fill_1 FILLER_9_45 ();
 sg13g2_fill_1 FILLER_9_51 ();
 sg13g2_fill_1 FILLER_9_57 ();
 sg13g2_fill_2 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_69 ();
 sg13g2_decap_8 FILLER_9_76 ();
 sg13g2_decap_8 FILLER_9_92 ();
 sg13g2_fill_2 FILLER_9_99 ();
 sg13g2_fill_1 FILLER_9_101 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_4 FILLER_9_137 ();
 sg13g2_fill_1 FILLER_9_141 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_fill_2 FILLER_9_161 ();
 sg13g2_fill_1 FILLER_9_163 ();
 sg13g2_fill_2 FILLER_9_174 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_4 FILLER_9_189 ();
 sg13g2_fill_2 FILLER_9_198 ();
 sg13g2_fill_2 FILLER_9_214 ();
 sg13g2_decap_8 FILLER_9_220 ();
 sg13g2_decap_4 FILLER_9_227 ();
 sg13g2_fill_1 FILLER_9_231 ();
 sg13g2_fill_2 FILLER_9_243 ();
 sg13g2_decap_8 FILLER_9_254 ();
 sg13g2_decap_8 FILLER_9_261 ();
 sg13g2_decap_4 FILLER_9_268 ();
 sg13g2_fill_1 FILLER_9_272 ();
 sg13g2_fill_1 FILLER_9_278 ();
 sg13g2_decap_8 FILLER_9_293 ();
 sg13g2_decap_4 FILLER_9_300 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_4 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_358 ();
 sg13g2_fill_2 FILLER_9_365 ();
 sg13g2_fill_1 FILLER_9_367 ();
 sg13g2_fill_2 FILLER_9_377 ();
 sg13g2_decap_8 FILLER_9_415 ();
 sg13g2_decap_8 FILLER_9_422 ();
 sg13g2_fill_2 FILLER_9_429 ();
 sg13g2_decap_8 FILLER_9_447 ();
 sg13g2_decap_8 FILLER_9_454 ();
 sg13g2_decap_4 FILLER_9_478 ();
 sg13g2_fill_2 FILLER_9_482 ();
 sg13g2_decap_8 FILLER_9_489 ();
 sg13g2_fill_2 FILLER_9_496 ();
 sg13g2_fill_1 FILLER_9_512 ();
 sg13g2_decap_8 FILLER_9_521 ();
 sg13g2_fill_1 FILLER_9_528 ();
 sg13g2_decap_8 FILLER_9_548 ();
 sg13g2_decap_4 FILLER_9_555 ();
 sg13g2_fill_1 FILLER_9_564 ();
 sg13g2_decap_8 FILLER_9_569 ();
 sg13g2_decap_8 FILLER_9_576 ();
 sg13g2_fill_2 FILLER_9_583 ();
 sg13g2_decap_4 FILLER_9_617 ();
 sg13g2_fill_1 FILLER_9_621 ();
 sg13g2_decap_4 FILLER_9_639 ();
 sg13g2_fill_1 FILLER_9_676 ();
 sg13g2_decap_8 FILLER_9_688 ();
 sg13g2_fill_2 FILLER_9_713 ();
 sg13g2_decap_8 FILLER_9_719 ();
 sg13g2_decap_4 FILLER_9_726 ();
 sg13g2_decap_4 FILLER_9_735 ();
 sg13g2_fill_1 FILLER_9_739 ();
 sg13g2_fill_2 FILLER_9_758 ();
 sg13g2_fill_1 FILLER_9_760 ();
 sg13g2_fill_1 FILLER_9_770 ();
 sg13g2_decap_8 FILLER_9_803 ();
 sg13g2_decap_4 FILLER_9_840 ();
 sg13g2_decap_8 FILLER_9_871 ();
 sg13g2_fill_2 FILLER_9_878 ();
 sg13g2_decap_8 FILLER_9_894 ();
 sg13g2_decap_4 FILLER_9_901 ();
 sg13g2_decap_4 FILLER_9_932 ();
 sg13g2_fill_2 FILLER_9_966 ();
 sg13g2_fill_2 FILLER_9_995 ();
 sg13g2_fill_2 FILLER_10_8 ();
 sg13g2_fill_1 FILLER_10_10 ();
 sg13g2_fill_2 FILLER_10_38 ();
 sg13g2_decap_8 FILLER_10_43 ();
 sg13g2_decap_8 FILLER_10_50 ();
 sg13g2_fill_1 FILLER_10_57 ();
 sg13g2_decap_8 FILLER_10_81 ();
 sg13g2_decap_8 FILLER_10_88 ();
 sg13g2_decap_8 FILLER_10_100 ();
 sg13g2_fill_2 FILLER_10_115 ();
 sg13g2_fill_1 FILLER_10_117 ();
 sg13g2_decap_8 FILLER_10_124 ();
 sg13g2_decap_8 FILLER_10_131 ();
 sg13g2_decap_4 FILLER_10_138 ();
 sg13g2_fill_1 FILLER_10_142 ();
 sg13g2_fill_2 FILLER_10_149 ();
 sg13g2_fill_1 FILLER_10_156 ();
 sg13g2_decap_8 FILLER_10_162 ();
 sg13g2_decap_4 FILLER_10_169 ();
 sg13g2_fill_1 FILLER_10_173 ();
 sg13g2_decap_4 FILLER_10_179 ();
 sg13g2_fill_2 FILLER_10_183 ();
 sg13g2_decap_8 FILLER_10_191 ();
 sg13g2_decap_8 FILLER_10_198 ();
 sg13g2_fill_2 FILLER_10_205 ();
 sg13g2_fill_1 FILLER_10_215 ();
 sg13g2_decap_8 FILLER_10_230 ();
 sg13g2_decap_4 FILLER_10_237 ();
 sg13g2_fill_2 FILLER_10_241 ();
 sg13g2_decap_8 FILLER_10_262 ();
 sg13g2_decap_8 FILLER_10_269 ();
 sg13g2_decap_8 FILLER_10_276 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_fill_2 FILLER_10_294 ();
 sg13g2_decap_4 FILLER_10_301 ();
 sg13g2_fill_1 FILLER_10_305 ();
 sg13g2_decap_8 FILLER_10_316 ();
 sg13g2_fill_2 FILLER_10_327 ();
 sg13g2_fill_1 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_349 ();
 sg13g2_fill_1 FILLER_10_356 ();
 sg13g2_fill_1 FILLER_10_367 ();
 sg13g2_fill_2 FILLER_10_380 ();
 sg13g2_fill_2 FILLER_10_393 ();
 sg13g2_decap_8 FILLER_10_416 ();
 sg13g2_fill_2 FILLER_10_423 ();
 sg13g2_decap_8 FILLER_10_446 ();
 sg13g2_decap_8 FILLER_10_480 ();
 sg13g2_decap_8 FILLER_10_487 ();
 sg13g2_decap_8 FILLER_10_494 ();
 sg13g2_decap_4 FILLER_10_501 ();
 sg13g2_fill_1 FILLER_10_510 ();
 sg13g2_fill_1 FILLER_10_545 ();
 sg13g2_decap_8 FILLER_10_558 ();
 sg13g2_decap_8 FILLER_10_565 ();
 sg13g2_decap_4 FILLER_10_572 ();
 sg13g2_decap_8 FILLER_10_583 ();
 sg13g2_decap_4 FILLER_10_590 ();
 sg13g2_fill_1 FILLER_10_594 ();
 sg13g2_decap_8 FILLER_10_599 ();
 sg13g2_decap_8 FILLER_10_606 ();
 sg13g2_fill_2 FILLER_10_613 ();
 sg13g2_fill_1 FILLER_10_615 ();
 sg13g2_fill_1 FILLER_10_643 ();
 sg13g2_fill_1 FILLER_10_685 ();
 sg13g2_fill_1 FILLER_10_743 ();
 sg13g2_fill_1 FILLER_10_771 ();
 sg13g2_fill_1 FILLER_10_777 ();
 sg13g2_fill_1 FILLER_10_781 ();
 sg13g2_fill_2 FILLER_10_786 ();
 sg13g2_fill_2 FILLER_10_801 ();
 sg13g2_fill_1 FILLER_10_803 ();
 sg13g2_decap_4 FILLER_10_836 ();
 sg13g2_fill_2 FILLER_10_840 ();
 sg13g2_fill_1 FILLER_10_847 ();
 sg13g2_decap_8 FILLER_10_861 ();
 sg13g2_decap_4 FILLER_10_901 ();
 sg13g2_fill_1 FILLER_10_905 ();
 sg13g2_fill_1 FILLER_10_940 ();
 sg13g2_fill_1 FILLER_10_950 ();
 sg13g2_decap_8 FILLER_10_960 ();
 sg13g2_decap_4 FILLER_10_967 ();
 sg13g2_fill_1 FILLER_10_971 ();
 sg13g2_decap_8 FILLER_10_985 ();
 sg13g2_fill_2 FILLER_10_992 ();
 sg13g2_decap_8 FILLER_10_1021 ();
 sg13g2_fill_1 FILLER_10_1028 ();
 sg13g2_fill_2 FILLER_11_4 ();
 sg13g2_fill_1 FILLER_11_6 ();
 sg13g2_decap_4 FILLER_11_17 ();
 sg13g2_fill_2 FILLER_11_29 ();
 sg13g2_decap_8 FILLER_11_41 ();
 sg13g2_fill_2 FILLER_11_48 ();
 sg13g2_decap_8 FILLER_11_54 ();
 sg13g2_decap_4 FILLER_11_61 ();
 sg13g2_fill_1 FILLER_11_65 ();
 sg13g2_decap_8 FILLER_11_71 ();
 sg13g2_decap_4 FILLER_11_78 ();
 sg13g2_fill_1 FILLER_11_82 ();
 sg13g2_decap_8 FILLER_11_94 ();
 sg13g2_decap_8 FILLER_11_101 ();
 sg13g2_decap_4 FILLER_11_108 ();
 sg13g2_decap_4 FILLER_11_122 ();
 sg13g2_fill_2 FILLER_11_126 ();
 sg13g2_decap_4 FILLER_11_137 ();
 sg13g2_fill_1 FILLER_11_141 ();
 sg13g2_fill_1 FILLER_11_148 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_4 FILLER_11_168 ();
 sg13g2_fill_1 FILLER_11_177 ();
 sg13g2_decap_8 FILLER_11_197 ();
 sg13g2_fill_1 FILLER_11_215 ();
 sg13g2_fill_2 FILLER_11_222 ();
 sg13g2_fill_1 FILLER_11_224 ();
 sg13g2_decap_4 FILLER_11_229 ();
 sg13g2_decap_4 FILLER_11_237 ();
 sg13g2_fill_2 FILLER_11_241 ();
 sg13g2_fill_2 FILLER_11_247 ();
 sg13g2_fill_1 FILLER_11_249 ();
 sg13g2_fill_2 FILLER_11_255 ();
 sg13g2_decap_4 FILLER_11_261 ();
 sg13g2_fill_2 FILLER_11_279 ();
 sg13g2_fill_1 FILLER_11_281 ();
 sg13g2_decap_8 FILLER_11_311 ();
 sg13g2_fill_1 FILLER_11_318 ();
 sg13g2_fill_1 FILLER_11_355 ();
 sg13g2_decap_4 FILLER_11_367 ();
 sg13g2_fill_1 FILLER_11_371 ();
 sg13g2_fill_2 FILLER_11_390 ();
 sg13g2_fill_1 FILLER_11_392 ();
 sg13g2_decap_4 FILLER_11_415 ();
 sg13g2_decap_8 FILLER_11_450 ();
 sg13g2_decap_8 FILLER_11_483 ();
 sg13g2_decap_4 FILLER_11_490 ();
 sg13g2_fill_1 FILLER_11_494 ();
 sg13g2_decap_8 FILLER_11_519 ();
 sg13g2_decap_8 FILLER_11_526 ();
 sg13g2_decap_4 FILLER_11_533 ();
 sg13g2_fill_1 FILLER_11_537 ();
 sg13g2_fill_2 FILLER_11_543 ();
 sg13g2_fill_1 FILLER_11_545 ();
 sg13g2_decap_8 FILLER_11_559 ();
 sg13g2_fill_1 FILLER_11_579 ();
 sg13g2_decap_8 FILLER_11_607 ();
 sg13g2_fill_1 FILLER_11_614 ();
 sg13g2_decap_8 FILLER_11_647 ();
 sg13g2_decap_8 FILLER_11_663 ();
 sg13g2_decap_4 FILLER_11_670 ();
 sg13g2_fill_2 FILLER_11_674 ();
 sg13g2_fill_1 FILLER_11_706 ();
 sg13g2_decap_4 FILLER_11_711 ();
 sg13g2_fill_2 FILLER_11_715 ();
 sg13g2_fill_2 FILLER_11_753 ();
 sg13g2_decap_4 FILLER_11_773 ();
 sg13g2_fill_2 FILLER_11_833 ();
 sg13g2_fill_1 FILLER_11_835 ();
 sg13g2_fill_1 FILLER_11_868 ();
 sg13g2_decap_4 FILLER_11_900 ();
 sg13g2_fill_2 FILLER_11_926 ();
 sg13g2_decap_8 FILLER_11_953 ();
 sg13g2_decap_4 FILLER_11_960 ();
 sg13g2_fill_1 FILLER_11_964 ();
 sg13g2_fill_2 FILLER_11_985 ();
 sg13g2_fill_1 FILLER_11_987 ();
 sg13g2_fill_2 FILLER_12_4 ();
 sg13g2_fill_1 FILLER_12_6 ();
 sg13g2_decap_4 FILLER_12_21 ();
 sg13g2_fill_1 FILLER_12_44 ();
 sg13g2_fill_2 FILLER_12_51 ();
 sg13g2_fill_1 FILLER_12_53 ();
 sg13g2_decap_8 FILLER_12_62 ();
 sg13g2_fill_2 FILLER_12_69 ();
 sg13g2_fill_1 FILLER_12_71 ();
 sg13g2_fill_2 FILLER_12_76 ();
 sg13g2_decap_8 FILLER_12_88 ();
 sg13g2_decap_8 FILLER_12_95 ();
 sg13g2_decap_8 FILLER_12_102 ();
 sg13g2_decap_8 FILLER_12_124 ();
 sg13g2_fill_2 FILLER_12_131 ();
 sg13g2_decap_8 FILLER_12_137 ();
 sg13g2_decap_4 FILLER_12_144 ();
 sg13g2_decap_8 FILLER_12_162 ();
 sg13g2_decap_8 FILLER_12_169 ();
 sg13g2_decap_4 FILLER_12_176 ();
 sg13g2_fill_1 FILLER_12_180 ();
 sg13g2_decap_8 FILLER_12_192 ();
 sg13g2_decap_8 FILLER_12_199 ();
 sg13g2_fill_1 FILLER_12_206 ();
 sg13g2_decap_8 FILLER_12_216 ();
 sg13g2_decap_8 FILLER_12_223 ();
 sg13g2_decap_4 FILLER_12_230 ();
 sg13g2_decap_8 FILLER_12_244 ();
 sg13g2_decap_8 FILLER_12_251 ();
 sg13g2_fill_2 FILLER_12_258 ();
 sg13g2_fill_1 FILLER_12_260 ();
 sg13g2_decap_8 FILLER_12_278 ();
 sg13g2_decap_8 FILLER_12_285 ();
 sg13g2_decap_8 FILLER_12_292 ();
 sg13g2_decap_8 FILLER_12_303 ();
 sg13g2_decap_8 FILLER_12_310 ();
 sg13g2_decap_8 FILLER_12_317 ();
 sg13g2_decap_8 FILLER_12_324 ();
 sg13g2_fill_2 FILLER_12_331 ();
 sg13g2_fill_1 FILLER_12_346 ();
 sg13g2_fill_2 FILLER_12_356 ();
 sg13g2_fill_1 FILLER_12_358 ();
 sg13g2_fill_2 FILLER_12_373 ();
 sg13g2_fill_1 FILLER_12_375 ();
 sg13g2_decap_8 FILLER_12_381 ();
 sg13g2_fill_2 FILLER_12_388 ();
 sg13g2_fill_1 FILLER_12_395 ();
 sg13g2_decap_8 FILLER_12_405 ();
 sg13g2_decap_8 FILLER_12_412 ();
 sg13g2_decap_8 FILLER_12_444 ();
 sg13g2_decap_8 FILLER_12_451 ();
 sg13g2_decap_4 FILLER_12_471 ();
 sg13g2_decap_8 FILLER_12_489 ();
 sg13g2_fill_2 FILLER_12_496 ();
 sg13g2_fill_1 FILLER_12_498 ();
 sg13g2_decap_8 FILLER_12_520 ();
 sg13g2_decap_8 FILLER_12_527 ();
 sg13g2_decap_8 FILLER_12_534 ();
 sg13g2_decap_8 FILLER_12_541 ();
 sg13g2_fill_2 FILLER_12_548 ();
 sg13g2_fill_1 FILLER_12_566 ();
 sg13g2_fill_1 FILLER_12_581 ();
 sg13g2_fill_1 FILLER_12_609 ();
 sg13g2_decap_8 FILLER_12_646 ();
 sg13g2_fill_1 FILLER_12_658 ();
 sg13g2_decap_4 FILLER_12_676 ();
 sg13g2_fill_2 FILLER_12_680 ();
 sg13g2_fill_2 FILLER_12_697 ();
 sg13g2_decap_8 FILLER_12_708 ();
 sg13g2_fill_1 FILLER_12_715 ();
 sg13g2_decap_4 FILLER_12_744 ();
 sg13g2_fill_2 FILLER_12_748 ();
 sg13g2_decap_4 FILLER_12_754 ();
 sg13g2_decap_8 FILLER_12_804 ();
 sg13g2_fill_1 FILLER_12_811 ();
 sg13g2_fill_2 FILLER_12_839 ();
 sg13g2_fill_2 FILLER_12_881 ();
 sg13g2_fill_1 FILLER_12_883 ();
 sg13g2_fill_1 FILLER_12_911 ();
 sg13g2_decap_8 FILLER_12_944 ();
 sg13g2_fill_2 FILLER_12_951 ();
 sg13g2_fill_1 FILLER_12_953 ();
 sg13g2_decap_8 FILLER_12_1021 ();
 sg13g2_fill_1 FILLER_12_1028 ();
 sg13g2_fill_2 FILLER_13_0 ();
 sg13g2_fill_1 FILLER_13_2 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_fill_2 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_46 ();
 sg13g2_decap_4 FILLER_13_59 ();
 sg13g2_fill_2 FILLER_13_63 ();
 sg13g2_decap_4 FILLER_13_82 ();
 sg13g2_fill_2 FILLER_13_95 ();
 sg13g2_decap_4 FILLER_13_101 ();
 sg13g2_fill_2 FILLER_13_105 ();
 sg13g2_decap_4 FILLER_13_138 ();
 sg13g2_fill_2 FILLER_13_142 ();
 sg13g2_fill_2 FILLER_13_167 ();
 sg13g2_fill_2 FILLER_13_173 ();
 sg13g2_fill_1 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_184 ();
 sg13g2_fill_1 FILLER_13_191 ();
 sg13g2_decap_8 FILLER_13_201 ();
 sg13g2_fill_2 FILLER_13_222 ();
 sg13g2_fill_1 FILLER_13_224 ();
 sg13g2_fill_2 FILLER_13_230 ();
 sg13g2_decap_4 FILLER_13_245 ();
 sg13g2_fill_2 FILLER_13_249 ();
 sg13g2_decap_4 FILLER_13_256 ();
 sg13g2_fill_1 FILLER_13_273 ();
 sg13g2_fill_1 FILLER_13_295 ();
 sg13g2_decap_4 FILLER_13_301 ();
 sg13g2_fill_2 FILLER_13_305 ();
 sg13g2_decap_8 FILLER_13_311 ();
 sg13g2_decap_8 FILLER_13_318 ();
 sg13g2_fill_1 FILLER_13_325 ();
 sg13g2_fill_1 FILLER_13_343 ();
 sg13g2_fill_2 FILLER_13_351 ();
 sg13g2_fill_1 FILLER_13_353 ();
 sg13g2_fill_2 FILLER_13_389 ();
 sg13g2_fill_1 FILLER_13_391 ();
 sg13g2_fill_2 FILLER_13_424 ();
 sg13g2_decap_4 FILLER_13_437 ();
 sg13g2_decap_8 FILLER_13_446 ();
 sg13g2_decap_4 FILLER_13_453 ();
 sg13g2_fill_2 FILLER_13_457 ();
 sg13g2_fill_2 FILLER_13_482 ();
 sg13g2_fill_1 FILLER_13_488 ();
 sg13g2_decap_8 FILLER_13_494 ();
 sg13g2_fill_2 FILLER_13_501 ();
 sg13g2_decap_8 FILLER_13_515 ();
 sg13g2_decap_8 FILLER_13_522 ();
 sg13g2_decap_4 FILLER_13_540 ();
 sg13g2_fill_1 FILLER_13_606 ();
 sg13g2_fill_1 FILLER_13_621 ();
 sg13g2_fill_2 FILLER_13_643 ();
 sg13g2_fill_2 FILLER_13_758 ();
 sg13g2_fill_1 FILLER_13_760 ();
 sg13g2_fill_1 FILLER_13_808 ();
 sg13g2_fill_2 FILLER_13_931 ();
 sg13g2_fill_2 FILLER_14_4 ();
 sg13g2_fill_1 FILLER_14_6 ();
 sg13g2_decap_8 FILLER_14_17 ();
 sg13g2_decap_8 FILLER_14_24 ();
 sg13g2_fill_2 FILLER_14_31 ();
 sg13g2_fill_1 FILLER_14_33 ();
 sg13g2_decap_8 FILLER_14_38 ();
 sg13g2_decap_8 FILLER_14_45 ();
 sg13g2_decap_8 FILLER_14_69 ();
 sg13g2_fill_2 FILLER_14_76 ();
 sg13g2_fill_1 FILLER_14_78 ();
 sg13g2_fill_2 FILLER_14_89 ();
 sg13g2_decap_8 FILLER_14_100 ();
 sg13g2_decap_8 FILLER_14_107 ();
 sg13g2_decap_8 FILLER_14_122 ();
 sg13g2_fill_1 FILLER_14_129 ();
 sg13g2_decap_4 FILLER_14_135 ();
 sg13g2_decap_8 FILLER_14_143 ();
 sg13g2_fill_2 FILLER_14_150 ();
 sg13g2_fill_1 FILLER_14_152 ();
 sg13g2_decap_8 FILLER_14_158 ();
 sg13g2_decap_8 FILLER_14_165 ();
 sg13g2_decap_8 FILLER_14_172 ();
 sg13g2_fill_2 FILLER_14_179 ();
 sg13g2_decap_8 FILLER_14_186 ();
 sg13g2_fill_2 FILLER_14_193 ();
 sg13g2_decap_8 FILLER_14_204 ();
 sg13g2_fill_2 FILLER_14_211 ();
 sg13g2_fill_1 FILLER_14_213 ();
 sg13g2_decap_8 FILLER_14_218 ();
 sg13g2_fill_1 FILLER_14_225 ();
 sg13g2_fill_2 FILLER_14_236 ();
 sg13g2_fill_1 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_4 FILLER_14_259 ();
 sg13g2_fill_2 FILLER_14_263 ();
 sg13g2_decap_8 FILLER_14_270 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_4 FILLER_14_294 ();
 sg13g2_fill_1 FILLER_14_298 ();
 sg13g2_decap_8 FILLER_14_389 ();
 sg13g2_decap_8 FILLER_14_396 ();
 sg13g2_decap_8 FILLER_14_403 ();
 sg13g2_decap_8 FILLER_14_410 ();
 sg13g2_fill_1 FILLER_14_417 ();
 sg13g2_fill_2 FILLER_14_431 ();
 sg13g2_decap_8 FILLER_14_450 ();
 sg13g2_decap_8 FILLER_14_457 ();
 sg13g2_fill_2 FILLER_14_464 ();
 sg13g2_fill_1 FILLER_14_466 ();
 sg13g2_decap_8 FILLER_14_471 ();
 sg13g2_decap_8 FILLER_14_478 ();
 sg13g2_fill_1 FILLER_14_485 ();
 sg13g2_decap_8 FILLER_14_519 ();
 sg13g2_decap_8 FILLER_14_542 ();
 sg13g2_decap_8 FILLER_14_549 ();
 sg13g2_decap_8 FILLER_14_556 ();
 sg13g2_fill_1 FILLER_14_563 ();
 sg13g2_decap_8 FILLER_14_604 ();
 sg13g2_decap_4 FILLER_14_611 ();
 sg13g2_fill_1 FILLER_14_615 ();
 sg13g2_fill_1 FILLER_14_649 ();
 sg13g2_decap_8 FILLER_14_654 ();
 sg13g2_fill_2 FILLER_14_661 ();
 sg13g2_decap_8 FILLER_14_669 ();
 sg13g2_decap_8 FILLER_14_680 ();
 sg13g2_fill_1 FILLER_14_687 ();
 sg13g2_fill_2 FILLER_14_711 ();
 sg13g2_decap_4 FILLER_14_722 ();
 sg13g2_fill_1 FILLER_14_726 ();
 sg13g2_fill_2 FILLER_14_800 ();
 sg13g2_fill_1 FILLER_14_838 ();
 sg13g2_fill_2 FILLER_14_848 ();
 sg13g2_fill_1 FILLER_14_949 ();
 sg13g2_fill_1 FILLER_14_964 ();
 sg13g2_fill_1 FILLER_14_992 ();
 sg13g2_fill_2 FILLER_15_4 ();
 sg13g2_fill_1 FILLER_15_6 ();
 sg13g2_decap_4 FILLER_15_18 ();
 sg13g2_fill_2 FILLER_15_22 ();
 sg13g2_fill_1 FILLER_15_33 ();
 sg13g2_decap_4 FILLER_15_47 ();
 sg13g2_fill_2 FILLER_15_51 ();
 sg13g2_decap_8 FILLER_15_71 ();
 sg13g2_decap_8 FILLER_15_78 ();
 sg13g2_decap_8 FILLER_15_85 ();
 sg13g2_fill_1 FILLER_15_92 ();
 sg13g2_decap_8 FILLER_15_97 ();
 sg13g2_decap_8 FILLER_15_104 ();
 sg13g2_decap_8 FILLER_15_111 ();
 sg13g2_fill_2 FILLER_15_122 ();
 sg13g2_decap_8 FILLER_15_137 ();
 sg13g2_decap_8 FILLER_15_144 ();
 sg13g2_fill_1 FILLER_15_151 ();
 sg13g2_decap_8 FILLER_15_164 ();
 sg13g2_decap_8 FILLER_15_171 ();
 sg13g2_fill_1 FILLER_15_178 ();
 sg13g2_decap_8 FILLER_15_184 ();
 sg13g2_decap_4 FILLER_15_191 ();
 sg13g2_fill_1 FILLER_15_195 ();
 sg13g2_decap_4 FILLER_15_201 ();
 sg13g2_decap_4 FILLER_15_213 ();
 sg13g2_decap_8 FILLER_15_221 ();
 sg13g2_fill_1 FILLER_15_228 ();
 sg13g2_fill_1 FILLER_15_234 ();
 sg13g2_fill_2 FILLER_15_239 ();
 sg13g2_fill_1 FILLER_15_241 ();
 sg13g2_fill_1 FILLER_15_260 ();
 sg13g2_decap_8 FILLER_15_265 ();
 sg13g2_fill_2 FILLER_15_272 ();
 sg13g2_fill_1 FILLER_15_274 ();
 sg13g2_decap_8 FILLER_15_288 ();
 sg13g2_decap_8 FILLER_15_295 ();
 sg13g2_fill_2 FILLER_15_302 ();
 sg13g2_fill_1 FILLER_15_304 ();
 sg13g2_fill_1 FILLER_15_309 ();
 sg13g2_decap_8 FILLER_15_314 ();
 sg13g2_decap_8 FILLER_15_321 ();
 sg13g2_fill_2 FILLER_15_328 ();
 sg13g2_fill_1 FILLER_15_330 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_4 FILLER_15_364 ();
 sg13g2_fill_1 FILLER_15_368 ();
 sg13g2_decap_4 FILLER_15_382 ();
 sg13g2_fill_1 FILLER_15_386 ();
 sg13g2_decap_4 FILLER_15_391 ();
 sg13g2_decap_8 FILLER_15_407 ();
 sg13g2_fill_1 FILLER_15_414 ();
 sg13g2_fill_1 FILLER_15_459 ();
 sg13g2_decap_8 FILLER_15_480 ();
 sg13g2_decap_8 FILLER_15_487 ();
 sg13g2_decap_8 FILLER_15_494 ();
 sg13g2_fill_2 FILLER_15_501 ();
 sg13g2_fill_1 FILLER_15_503 ();
 sg13g2_decap_8 FILLER_15_513 ();
 sg13g2_decap_8 FILLER_15_520 ();
 sg13g2_fill_2 FILLER_15_527 ();
 sg13g2_fill_1 FILLER_15_534 ();
 sg13g2_decap_8 FILLER_15_562 ();
 sg13g2_decap_8 FILLER_15_569 ();
 sg13g2_decap_8 FILLER_15_576 ();
 sg13g2_fill_2 FILLER_15_583 ();
 sg13g2_fill_1 FILLER_15_585 ();
 sg13g2_decap_4 FILLER_15_617 ();
 sg13g2_fill_2 FILLER_15_625 ();
 sg13g2_fill_1 FILLER_15_627 ();
 sg13g2_decap_8 FILLER_15_633 ();
 sg13g2_fill_2 FILLER_15_640 ();
 sg13g2_fill_1 FILLER_15_642 ();
 sg13g2_decap_8 FILLER_15_662 ();
 sg13g2_decap_4 FILLER_15_669 ();
 sg13g2_fill_1 FILLER_15_673 ();
 sg13g2_fill_2 FILLER_15_692 ();
 sg13g2_fill_1 FILLER_15_694 ();
 sg13g2_fill_2 FILLER_15_722 ();
 sg13g2_fill_1 FILLER_15_724 ();
 sg13g2_fill_2 FILLER_15_730 ();
 sg13g2_fill_1 FILLER_15_732 ();
 sg13g2_fill_2 FILLER_15_739 ();
 sg13g2_fill_2 FILLER_15_768 ();
 sg13g2_fill_1 FILLER_15_770 ();
 sg13g2_fill_1 FILLER_15_784 ();
 sg13g2_fill_2 FILLER_15_794 ();
 sg13g2_fill_1 FILLER_15_805 ();
 sg13g2_fill_2 FILLER_15_824 ();
 sg13g2_decap_4 FILLER_15_867 ();
 sg13g2_fill_2 FILLER_15_871 ();
 sg13g2_fill_1 FILLER_15_926 ();
 sg13g2_fill_2 FILLER_15_951 ();
 sg13g2_fill_2 FILLER_15_980 ();
 sg13g2_fill_2 FILLER_15_1017 ();
 sg13g2_fill_1 FILLER_15_1019 ();
 sg13g2_fill_2 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_2 ();
 sg13g2_decap_4 FILLER_16_43 ();
 sg13g2_fill_2 FILLER_16_69 ();
 sg13g2_fill_2 FILLER_16_79 ();
 sg13g2_fill_1 FILLER_16_81 ();
 sg13g2_decap_8 FILLER_16_102 ();
 sg13g2_fill_1 FILLER_16_109 ();
 sg13g2_fill_1 FILLER_16_119 ();
 sg13g2_decap_4 FILLER_16_138 ();
 sg13g2_fill_2 FILLER_16_142 ();
 sg13g2_fill_2 FILLER_16_168 ();
 sg13g2_fill_1 FILLER_16_170 ();
 sg13g2_fill_2 FILLER_16_197 ();
 sg13g2_decap_8 FILLER_16_204 ();
 sg13g2_fill_2 FILLER_16_211 ();
 sg13g2_decap_8 FILLER_16_218 ();
 sg13g2_decap_8 FILLER_16_225 ();
 sg13g2_decap_4 FILLER_16_240 ();
 sg13g2_fill_1 FILLER_16_244 ();
 sg13g2_fill_2 FILLER_16_260 ();
 sg13g2_fill_2 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_275 ();
 sg13g2_fill_1 FILLER_16_287 ();
 sg13g2_fill_2 FILLER_16_297 ();
 sg13g2_fill_1 FILLER_16_299 ();
 sg13g2_fill_1 FILLER_16_304 ();
 sg13g2_decap_4 FILLER_16_345 ();
 sg13g2_fill_2 FILLER_16_361 ();
 sg13g2_fill_1 FILLER_16_363 ();
 sg13g2_fill_2 FILLER_16_371 ();
 sg13g2_fill_1 FILLER_16_373 ();
 sg13g2_decap_4 FILLER_16_383 ();
 sg13g2_fill_1 FILLER_16_419 ();
 sg13g2_fill_2 FILLER_16_460 ();
 sg13g2_fill_1 FILLER_16_462 ();
 sg13g2_decap_8 FILLER_16_504 ();
 sg13g2_decap_4 FILLER_16_511 ();
 sg13g2_fill_1 FILLER_16_520 ();
 sg13g2_fill_2 FILLER_16_526 ();
 sg13g2_decap_4 FILLER_16_546 ();
 sg13g2_decap_8 FILLER_16_571 ();
 sg13g2_fill_1 FILLER_16_578 ();
 sg13g2_fill_1 FILLER_16_582 ();
 sg13g2_fill_2 FILLER_16_587 ();
 sg13g2_fill_1 FILLER_16_589 ();
 sg13g2_decap_4 FILLER_16_630 ();
 sg13g2_fill_2 FILLER_16_754 ();
 sg13g2_fill_1 FILLER_16_756 ();
 sg13g2_decap_4 FILLER_16_761 ();
 sg13g2_fill_2 FILLER_16_819 ();
 sg13g2_fill_1 FILLER_16_821 ();
 sg13g2_fill_2 FILLER_16_827 ();
 sg13g2_fill_1 FILLER_16_829 ();
 sg13g2_decap_8 FILLER_16_835 ();
 sg13g2_decap_8 FILLER_16_842 ();
 sg13g2_fill_2 FILLER_16_849 ();
 sg13g2_fill_1 FILLER_16_851 ();
 sg13g2_fill_1 FILLER_16_860 ();
 sg13g2_decap_4 FILLER_16_865 ();
 sg13g2_fill_2 FILLER_16_869 ();
 sg13g2_decap_4 FILLER_16_892 ();
 sg13g2_fill_2 FILLER_16_926 ();
 sg13g2_fill_1 FILLER_16_973 ();
 sg13g2_fill_1 FILLER_16_988 ();
 sg13g2_decap_8 FILLER_16_1021 ();
 sg13g2_fill_1 FILLER_16_1028 ();
 sg13g2_fill_2 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_2 ();
 sg13g2_fill_2 FILLER_17_27 ();
 sg13g2_decap_8 FILLER_17_44 ();
 sg13g2_decap_8 FILLER_17_51 ();
 sg13g2_fill_2 FILLER_17_63 ();
 sg13g2_fill_2 FILLER_17_73 ();
 sg13g2_fill_1 FILLER_17_75 ();
 sg13g2_decap_8 FILLER_17_116 ();
 sg13g2_decap_4 FILLER_17_123 ();
 sg13g2_fill_1 FILLER_17_127 ();
 sg13g2_decap_8 FILLER_17_132 ();
 sg13g2_decap_4 FILLER_17_139 ();
 sg13g2_fill_2 FILLER_17_143 ();
 sg13g2_decap_8 FILLER_17_170 ();
 sg13g2_decap_8 FILLER_17_177 ();
 sg13g2_fill_2 FILLER_17_184 ();
 sg13g2_fill_1 FILLER_17_186 ();
 sg13g2_fill_2 FILLER_17_210 ();
 sg13g2_fill_1 FILLER_17_212 ();
 sg13g2_decap_8 FILLER_17_249 ();
 sg13g2_decap_8 FILLER_17_256 ();
 sg13g2_decap_8 FILLER_17_263 ();
 sg13g2_fill_1 FILLER_17_270 ();
 sg13g2_decap_4 FILLER_17_275 ();
 sg13g2_fill_1 FILLER_17_279 ();
 sg13g2_decap_8 FILLER_17_304 ();
 sg13g2_decap_4 FILLER_17_311 ();
 sg13g2_fill_2 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_328 ();
 sg13g2_decap_8 FILLER_17_335 ();
 sg13g2_fill_2 FILLER_17_342 ();
 sg13g2_fill_1 FILLER_17_344 ();
 sg13g2_fill_2 FILLER_17_354 ();
 sg13g2_fill_1 FILLER_17_356 ();
 sg13g2_fill_2 FILLER_17_361 ();
 sg13g2_decap_8 FILLER_17_390 ();
 sg13g2_decap_4 FILLER_17_397 ();
 sg13g2_decap_8 FILLER_17_408 ();
 sg13g2_fill_2 FILLER_17_415 ();
 sg13g2_decap_8 FILLER_17_422 ();
 sg13g2_fill_1 FILLER_17_429 ();
 sg13g2_fill_2 FILLER_17_451 ();
 sg13g2_decap_8 FILLER_17_461 ();
 sg13g2_fill_2 FILLER_17_468 ();
 sg13g2_decap_8 FILLER_17_478 ();
 sg13g2_decap_4 FILLER_17_485 ();
 sg13g2_fill_2 FILLER_17_520 ();
 sg13g2_decap_8 FILLER_17_526 ();
 sg13g2_fill_2 FILLER_17_538 ();
 sg13g2_fill_1 FILLER_17_540 ();
 sg13g2_fill_2 FILLER_17_546 ();
 sg13g2_fill_1 FILLER_17_555 ();
 sg13g2_fill_2 FILLER_17_615 ();
 sg13g2_fill_1 FILLER_17_617 ();
 sg13g2_fill_1 FILLER_17_645 ();
 sg13g2_decap_4 FILLER_17_668 ();
 sg13g2_fill_2 FILLER_17_677 ();
 sg13g2_fill_1 FILLER_17_684 ();
 sg13g2_fill_2 FILLER_17_690 ();
 sg13g2_fill_1 FILLER_17_716 ();
 sg13g2_fill_1 FILLER_17_722 ();
 sg13g2_fill_2 FILLER_17_773 ();
 sg13g2_fill_1 FILLER_17_780 ();
 sg13g2_decap_8 FILLER_17_786 ();
 sg13g2_decap_8 FILLER_17_828 ();
 sg13g2_fill_1 FILLER_17_835 ();
 sg13g2_decap_4 FILLER_17_841 ();
 sg13g2_fill_2 FILLER_17_845 ();
 sg13g2_decap_4 FILLER_17_919 ();
 sg13g2_fill_1 FILLER_17_941 ();
 sg13g2_fill_2 FILLER_17_1000 ();
 sg13g2_fill_2 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_2 ();
 sg13g2_fill_1 FILLER_18_48 ();
 sg13g2_decap_8 FILLER_18_76 ();
 sg13g2_decap_8 FILLER_18_83 ();
 sg13g2_decap_8 FILLER_18_90 ();
 sg13g2_fill_2 FILLER_18_97 ();
 sg13g2_fill_1 FILLER_18_102 ();
 sg13g2_fill_2 FILLER_18_109 ();
 sg13g2_fill_1 FILLER_18_111 ();
 sg13g2_decap_8 FILLER_18_116 ();
 sg13g2_fill_2 FILLER_18_123 ();
 sg13g2_fill_1 FILLER_18_125 ();
 sg13g2_decap_8 FILLER_18_136 ();
 sg13g2_decap_8 FILLER_18_143 ();
 sg13g2_decap_8 FILLER_18_150 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_fill_1 FILLER_18_182 ();
 sg13g2_fill_2 FILLER_18_195 ();
 sg13g2_fill_1 FILLER_18_205 ();
 sg13g2_decap_8 FILLER_18_211 ();
 sg13g2_decap_8 FILLER_18_218 ();
 sg13g2_fill_2 FILLER_18_225 ();
 sg13g2_decap_4 FILLER_18_231 ();
 sg13g2_fill_1 FILLER_18_235 ();
 sg13g2_decap_8 FILLER_18_267 ();
 sg13g2_decap_8 FILLER_18_274 ();
 sg13g2_decap_8 FILLER_18_281 ();
 sg13g2_decap_8 FILLER_18_299 ();
 sg13g2_decap_8 FILLER_18_306 ();
 sg13g2_decap_4 FILLER_18_313 ();
 sg13g2_decap_8 FILLER_18_327 ();
 sg13g2_decap_8 FILLER_18_334 ();
 sg13g2_decap_8 FILLER_18_341 ();
 sg13g2_decap_4 FILLER_18_348 ();
 sg13g2_fill_2 FILLER_18_356 ();
 sg13g2_fill_1 FILLER_18_358 ();
 sg13g2_fill_1 FILLER_18_364 ();
 sg13g2_fill_2 FILLER_18_375 ();
 sg13g2_fill_1 FILLER_18_377 ();
 sg13g2_decap_8 FILLER_18_387 ();
 sg13g2_decap_8 FILLER_18_394 ();
 sg13g2_fill_2 FILLER_18_401 ();
 sg13g2_fill_1 FILLER_18_403 ();
 sg13g2_fill_1 FILLER_18_431 ();
 sg13g2_fill_1 FILLER_18_452 ();
 sg13g2_decap_8 FILLER_18_461 ();
 sg13g2_decap_8 FILLER_18_531 ();
 sg13g2_fill_2 FILLER_18_538 ();
 sg13g2_fill_1 FILLER_18_540 ();
 sg13g2_fill_2 FILLER_18_579 ();
 sg13g2_fill_1 FILLER_18_600 ();
 sg13g2_decap_4 FILLER_18_614 ();
 sg13g2_fill_1 FILLER_18_637 ();
 sg13g2_fill_2 FILLER_18_674 ();
 sg13g2_fill_2 FILLER_18_695 ();
 sg13g2_fill_1 FILLER_18_732 ();
 sg13g2_fill_1 FILLER_18_762 ();
 sg13g2_decap_8 FILLER_18_785 ();
 sg13g2_decap_8 FILLER_18_792 ();
 sg13g2_fill_2 FILLER_18_799 ();
 sg13g2_fill_1 FILLER_18_801 ();
 sg13g2_fill_2 FILLER_18_813 ();
 sg13g2_decap_4 FILLER_18_819 ();
 sg13g2_fill_1 FILLER_18_823 ();
 sg13g2_fill_2 FILLER_18_831 ();
 sg13g2_fill_2 FILLER_18_842 ();
 sg13g2_fill_1 FILLER_18_844 ();
 sg13g2_fill_2 FILLER_18_849 ();
 sg13g2_decap_4 FILLER_18_875 ();
 sg13g2_fill_1 FILLER_18_879 ();
 sg13g2_fill_1 FILLER_18_903 ();
 sg13g2_fill_2 FILLER_18_908 ();
 sg13g2_decap_4 FILLER_18_915 ();
 sg13g2_fill_1 FILLER_18_919 ();
 sg13g2_fill_2 FILLER_18_925 ();
 sg13g2_decap_8 FILLER_18_959 ();
 sg13g2_fill_2 FILLER_18_966 ();
 sg13g2_fill_1 FILLER_18_968 ();
 sg13g2_fill_2 FILLER_18_977 ();
 sg13g2_fill_2 FILLER_18_983 ();
 sg13g2_fill_1 FILLER_18_998 ();
 sg13g2_fill_2 FILLER_18_1013 ();
 sg13g2_fill_1 FILLER_18_1015 ();
 sg13g2_fill_2 FILLER_19_8 ();
 sg13g2_fill_1 FILLER_19_10 ();
 sg13g2_fill_2 FILLER_19_46 ();
 sg13g2_fill_1 FILLER_19_48 ();
 sg13g2_decap_8 FILLER_19_52 ();
 sg13g2_decap_4 FILLER_19_70 ();
 sg13g2_fill_2 FILLER_19_74 ();
 sg13g2_fill_1 FILLER_19_103 ();
 sg13g2_decap_4 FILLER_19_158 ();
 sg13g2_fill_1 FILLER_19_162 ();
 sg13g2_fill_2 FILLER_19_187 ();
 sg13g2_fill_1 FILLER_19_189 ();
 sg13g2_decap_4 FILLER_19_213 ();
 sg13g2_decap_8 FILLER_19_235 ();
 sg13g2_decap_4 FILLER_19_242 ();
 sg13g2_fill_1 FILLER_19_246 ();
 sg13g2_fill_1 FILLER_19_279 ();
 sg13g2_fill_2 FILLER_19_337 ();
 sg13g2_decap_8 FILLER_19_349 ();
 sg13g2_decap_4 FILLER_19_356 ();
 sg13g2_fill_2 FILLER_19_360 ();
 sg13g2_decap_8 FILLER_19_423 ();
 sg13g2_fill_1 FILLER_19_430 ();
 sg13g2_decap_4 FILLER_19_465 ();
 sg13g2_fill_1 FILLER_19_469 ();
 sg13g2_fill_2 FILLER_19_501 ();
 sg13g2_fill_2 FILLER_19_512 ();
 sg13g2_fill_1 FILLER_19_514 ();
 sg13g2_decap_8 FILLER_19_599 ();
 sg13g2_decap_4 FILLER_19_606 ();
 sg13g2_fill_1 FILLER_19_610 ();
 sg13g2_decap_4 FILLER_19_616 ();
 sg13g2_fill_2 FILLER_19_647 ();
 sg13g2_fill_1 FILLER_19_689 ();
 sg13g2_fill_1 FILLER_19_735 ();
 sg13g2_fill_2 FILLER_19_750 ();
 sg13g2_fill_2 FILLER_19_756 ();
 sg13g2_fill_1 FILLER_19_767 ();
 sg13g2_fill_2 FILLER_19_801 ();
 sg13g2_fill_2 FILLER_19_808 ();
 sg13g2_fill_1 FILLER_19_818 ();
 sg13g2_decap_8 FILLER_19_839 ();
 sg13g2_fill_2 FILLER_19_846 ();
 sg13g2_decap_8 FILLER_19_867 ();
 sg13g2_fill_2 FILLER_19_874 ();
 sg13g2_decap_4 FILLER_19_880 ();
 sg13g2_fill_1 FILLER_19_884 ();
 sg13g2_fill_2 FILLER_19_895 ();
 sg13g2_decap_8 FILLER_19_902 ();
 sg13g2_decap_4 FILLER_19_909 ();
 sg13g2_fill_1 FILLER_19_913 ();
 sg13g2_decap_8 FILLER_19_941 ();
 sg13g2_fill_2 FILLER_19_948 ();
 sg13g2_decap_8 FILLER_19_956 ();
 sg13g2_fill_2 FILLER_19_963 ();
 sg13g2_fill_1 FILLER_19_965 ();
 sg13g2_fill_1 FILLER_19_976 ();
 sg13g2_fill_2 FILLER_19_982 ();
 sg13g2_fill_2 FILLER_19_997 ();
 sg13g2_fill_2 FILLER_20_4 ();
 sg13g2_fill_1 FILLER_20_6 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_fill_2 FILLER_20_35 ();
 sg13g2_fill_2 FILLER_20_68 ();
 sg13g2_fill_2 FILLER_20_88 ();
 sg13g2_decap_4 FILLER_20_129 ();
 sg13g2_fill_2 FILLER_20_133 ();
 sg13g2_fill_2 FILLER_20_147 ();
 sg13g2_fill_1 FILLER_20_149 ();
 sg13g2_fill_1 FILLER_20_162 ();
 sg13g2_fill_2 FILLER_20_175 ();
 sg13g2_fill_2 FILLER_20_181 ();
 sg13g2_decap_8 FILLER_20_191 ();
 sg13g2_fill_2 FILLER_20_198 ();
 sg13g2_decap_8 FILLER_20_209 ();
 sg13g2_fill_1 FILLER_20_216 ();
 sg13g2_decap_8 FILLER_20_257 ();
 sg13g2_decap_8 FILLER_20_264 ();
 sg13g2_fill_2 FILLER_20_285 ();
 sg13g2_fill_2 FILLER_20_291 ();
 sg13g2_decap_8 FILLER_20_299 ();
 sg13g2_decap_4 FILLER_20_306 ();
 sg13g2_fill_2 FILLER_20_346 ();
 sg13g2_fill_1 FILLER_20_348 ();
 sg13g2_fill_1 FILLER_20_376 ();
 sg13g2_fill_2 FILLER_20_381 ();
 sg13g2_fill_2 FILLER_20_395 ();
 sg13g2_fill_1 FILLER_20_397 ();
 sg13g2_decap_8 FILLER_20_429 ();
 sg13g2_fill_1 FILLER_20_436 ();
 sg13g2_fill_1 FILLER_20_470 ();
 sg13g2_fill_1 FILLER_20_498 ();
 sg13g2_fill_2 FILLER_20_524 ();
 sg13g2_fill_2 FILLER_20_531 ();
 sg13g2_decap_4 FILLER_20_551 ();
 sg13g2_fill_2 FILLER_20_555 ();
 sg13g2_fill_2 FILLER_20_629 ();
 sg13g2_fill_1 FILLER_20_631 ();
 sg13g2_decap_8 FILLER_20_635 ();
 sg13g2_fill_1 FILLER_20_642 ();
 sg13g2_fill_2 FILLER_20_653 ();
 sg13g2_fill_2 FILLER_20_682 ();
 sg13g2_fill_1 FILLER_20_705 ();
 sg13g2_fill_1 FILLER_20_847 ();
 sg13g2_fill_2 FILLER_20_910 ();
 sg13g2_decap_4 FILLER_20_939 ();
 sg13g2_fill_1 FILLER_20_943 ();
 sg13g2_decap_8 FILLER_20_1019 ();
 sg13g2_fill_2 FILLER_20_1026 ();
 sg13g2_fill_1 FILLER_20_1028 ();
 sg13g2_fill_2 FILLER_21_4 ();
 sg13g2_fill_1 FILLER_21_6 ();
 sg13g2_decap_4 FILLER_21_21 ();
 sg13g2_fill_2 FILLER_21_25 ();
 sg13g2_fill_2 FILLER_21_38 ();
 sg13g2_fill_1 FILLER_21_70 ();
 sg13g2_fill_2 FILLER_21_79 ();
 sg13g2_fill_1 FILLER_21_121 ();
 sg13g2_fill_2 FILLER_21_155 ();
 sg13g2_fill_1 FILLER_21_188 ();
 sg13g2_decap_8 FILLER_21_197 ();
 sg13g2_decap_8 FILLER_21_208 ();
 sg13g2_decap_8 FILLER_21_215 ();
 sg13g2_fill_2 FILLER_21_222 ();
 sg13g2_fill_1 FILLER_21_224 ();
 sg13g2_decap_4 FILLER_21_230 ();
 sg13g2_fill_1 FILLER_21_234 ();
 sg13g2_fill_1 FILLER_21_272 ();
 sg13g2_decap_8 FILLER_21_297 ();
 sg13g2_decap_8 FILLER_21_304 ();
 sg13g2_decap_8 FILLER_21_311 ();
 sg13g2_fill_2 FILLER_21_318 ();
 sg13g2_fill_1 FILLER_21_320 ();
 sg13g2_fill_2 FILLER_21_326 ();
 sg13g2_fill_2 FILLER_21_333 ();
 sg13g2_fill_1 FILLER_21_335 ();
 sg13g2_decap_4 FILLER_21_344 ();
 sg13g2_fill_1 FILLER_21_348 ();
 sg13g2_fill_2 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_368 ();
 sg13g2_decap_4 FILLER_21_375 ();
 sg13g2_fill_1 FILLER_21_379 ();
 sg13g2_fill_2 FILLER_21_388 ();
 sg13g2_decap_8 FILLER_21_394 ();
 sg13g2_decap_4 FILLER_21_414 ();
 sg13g2_fill_1 FILLER_21_487 ();
 sg13g2_fill_1 FILLER_21_528 ();
 sg13g2_decap_8 FILLER_21_542 ();
 sg13g2_decap_4 FILLER_21_549 ();
 sg13g2_fill_2 FILLER_21_553 ();
 sg13g2_fill_1 FILLER_21_608 ();
 sg13g2_fill_2 FILLER_21_626 ();
 sg13g2_fill_1 FILLER_21_635 ();
 sg13g2_fill_2 FILLER_21_667 ();
 sg13g2_fill_2 FILLER_21_674 ();
 sg13g2_fill_2 FILLER_21_687 ();
 sg13g2_fill_1 FILLER_21_716 ();
 sg13g2_decap_8 FILLER_21_755 ();
 sg13g2_decap_8 FILLER_21_762 ();
 sg13g2_fill_2 FILLER_21_769 ();
 sg13g2_fill_1 FILLER_21_771 ();
 sg13g2_fill_1 FILLER_21_790 ();
 sg13g2_fill_2 FILLER_21_801 ();
 sg13g2_fill_2 FILLER_21_824 ();
 sg13g2_fill_2 FILLER_21_875 ();
 sg13g2_fill_1 FILLER_21_877 ();
 sg13g2_fill_2 FILLER_21_897 ();
 sg13g2_decap_4 FILLER_21_925 ();
 sg13g2_fill_2 FILLER_21_956 ();
 sg13g2_fill_1 FILLER_21_958 ();
 sg13g2_fill_2 FILLER_21_991 ();
 sg13g2_decap_8 FILLER_21_1021 ();
 sg13g2_fill_1 FILLER_21_1028 ();
 sg13g2_fill_2 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_2 ();
 sg13g2_fill_2 FILLER_22_17 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_fill_2 FILLER_22_42 ();
 sg13g2_fill_1 FILLER_22_53 ();
 sg13g2_fill_2 FILLER_22_60 ();
 sg13g2_fill_1 FILLER_22_62 ();
 sg13g2_decap_4 FILLER_22_72 ();
 sg13g2_fill_1 FILLER_22_76 ();
 sg13g2_decap_8 FILLER_22_88 ();
 sg13g2_decap_8 FILLER_22_95 ();
 sg13g2_decap_4 FILLER_22_102 ();
 sg13g2_fill_1 FILLER_22_106 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_4 FILLER_22_138 ();
 sg13g2_fill_1 FILLER_22_142 ();
 sg13g2_fill_2 FILLER_22_183 ();
 sg13g2_fill_1 FILLER_22_190 ();
 sg13g2_fill_2 FILLER_22_205 ();
 sg13g2_fill_1 FILLER_22_207 ();
 sg13g2_decap_4 FILLER_22_213 ();
 sg13g2_fill_1 FILLER_22_217 ();
 sg13g2_fill_2 FILLER_22_223 ();
 sg13g2_fill_2 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_249 ();
 sg13g2_decap_8 FILLER_22_256 ();
 sg13g2_decap_8 FILLER_22_263 ();
 sg13g2_fill_1 FILLER_22_270 ();
 sg13g2_fill_1 FILLER_22_300 ();
 sg13g2_fill_1 FILLER_22_318 ();
 sg13g2_decap_4 FILLER_22_345 ();
 sg13g2_decap_8 FILLER_22_355 ();
 sg13g2_decap_4 FILLER_22_362 ();
 sg13g2_fill_2 FILLER_22_366 ();
 sg13g2_fill_2 FILLER_22_372 ();
 sg13g2_fill_1 FILLER_22_374 ();
 sg13g2_decap_4 FILLER_22_408 ();
 sg13g2_fill_1 FILLER_22_412 ();
 sg13g2_decap_4 FILLER_22_431 ();
 sg13g2_fill_2 FILLER_22_435 ();
 sg13g2_fill_2 FILLER_22_449 ();
 sg13g2_fill_2 FILLER_22_488 ();
 sg13g2_fill_2 FILLER_22_517 ();
 sg13g2_fill_1 FILLER_22_519 ();
 sg13g2_decap_4 FILLER_22_549 ();
 sg13g2_fill_2 FILLER_22_553 ();
 sg13g2_fill_1 FILLER_22_563 ();
 sg13g2_decap_4 FILLER_22_650 ();
 sg13g2_fill_1 FILLER_22_654 ();
 sg13g2_fill_2 FILLER_22_713 ();
 sg13g2_fill_1 FILLER_22_742 ();
 sg13g2_decap_4 FILLER_22_758 ();
 sg13g2_fill_2 FILLER_22_762 ();
 sg13g2_fill_1 FILLER_22_800 ();
 sg13g2_fill_1 FILLER_22_809 ();
 sg13g2_decap_4 FILLER_22_846 ();
 sg13g2_fill_1 FILLER_22_859 ();
 sg13g2_decap_4 FILLER_22_868 ();
 sg13g2_fill_2 FILLER_22_876 ();
 sg13g2_fill_1 FILLER_22_878 ();
 sg13g2_fill_2 FILLER_22_933 ();
 sg13g2_fill_2 FILLER_22_960 ();
 sg13g2_fill_1 FILLER_22_962 ();
 sg13g2_fill_1 FILLER_22_989 ();
 sg13g2_decap_4 FILLER_22_993 ();
 sg13g2_fill_2 FILLER_23_8 ();
 sg13g2_fill_1 FILLER_23_10 ();
 sg13g2_decap_4 FILLER_23_15 ();
 sg13g2_fill_2 FILLER_23_19 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_4 FILLER_23_35 ();
 sg13g2_fill_1 FILLER_23_39 ();
 sg13g2_fill_1 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_100 ();
 sg13g2_fill_1 FILLER_23_107 ();
 sg13g2_fill_2 FILLER_23_113 ();
 sg13g2_fill_1 FILLER_23_115 ();
 sg13g2_decap_8 FILLER_23_124 ();
 sg13g2_decap_8 FILLER_23_131 ();
 sg13g2_fill_2 FILLER_23_145 ();
 sg13g2_fill_2 FILLER_23_181 ();
 sg13g2_fill_2 FILLER_23_195 ();
 sg13g2_fill_1 FILLER_23_197 ();
 sg13g2_decap_8 FILLER_23_226 ();
 sg13g2_fill_2 FILLER_23_233 ();
 sg13g2_fill_1 FILLER_23_235 ();
 sg13g2_decap_8 FILLER_23_244 ();
 sg13g2_fill_2 FILLER_23_251 ();
 sg13g2_fill_1 FILLER_23_253 ();
 sg13g2_fill_1 FILLER_23_260 ();
 sg13g2_decap_8 FILLER_23_267 ();
 sg13g2_fill_2 FILLER_23_274 ();
 sg13g2_decap_4 FILLER_23_297 ();
 sg13g2_fill_1 FILLER_23_307 ();
 sg13g2_fill_1 FILLER_23_318 ();
 sg13g2_decap_8 FILLER_23_323 ();
 sg13g2_fill_2 FILLER_23_342 ();
 sg13g2_fill_1 FILLER_23_344 ();
 sg13g2_decap_8 FILLER_23_363 ();
 sg13g2_decap_8 FILLER_23_370 ();
 sg13g2_decap_8 FILLER_23_377 ();
 sg13g2_fill_1 FILLER_23_384 ();
 sg13g2_fill_2 FILLER_23_412 ();
 sg13g2_decap_4 FILLER_23_429 ();
 sg13g2_fill_1 FILLER_23_433 ();
 sg13g2_fill_2 FILLER_23_446 ();
 sg13g2_fill_1 FILLER_23_448 ();
 sg13g2_decap_8 FILLER_23_459 ();
 sg13g2_fill_2 FILLER_23_466 ();
 sg13g2_fill_1 FILLER_23_468 ();
 sg13g2_decap_8 FILLER_23_478 ();
 sg13g2_fill_1 FILLER_23_499 ();
 sg13g2_decap_8 FILLER_23_504 ();
 sg13g2_fill_1 FILLER_23_511 ();
 sg13g2_decap_4 FILLER_23_527 ();
 sg13g2_decap_4 FILLER_23_555 ();
 sg13g2_fill_1 FILLER_23_559 ();
 sg13g2_fill_1 FILLER_23_594 ();
 sg13g2_decap_8 FILLER_23_605 ();
 sg13g2_fill_2 FILLER_23_612 ();
 sg13g2_fill_1 FILLER_23_655 ();
 sg13g2_fill_1 FILLER_23_667 ();
 sg13g2_decap_8 FILLER_23_673 ();
 sg13g2_fill_1 FILLER_23_680 ();
 sg13g2_fill_2 FILLER_23_701 ();
 sg13g2_fill_1 FILLER_23_703 ();
 sg13g2_decap_8 FILLER_23_712 ();
 sg13g2_fill_2 FILLER_23_731 ();
 sg13g2_fill_1 FILLER_23_733 ();
 sg13g2_decap_4 FILLER_23_765 ();
 sg13g2_decap_4 FILLER_23_773 ();
 sg13g2_decap_8 FILLER_23_791 ();
 sg13g2_decap_4 FILLER_23_798 ();
 sg13g2_fill_1 FILLER_23_802 ();
 sg13g2_fill_1 FILLER_23_830 ();
 sg13g2_decap_4 FILLER_23_835 ();
 sg13g2_fill_2 FILLER_23_842 ();
 sg13g2_fill_1 FILLER_23_844 ();
 sg13g2_fill_2 FILLER_23_895 ();
 sg13g2_fill_1 FILLER_23_910 ();
 sg13g2_fill_2 FILLER_23_934 ();
 sg13g2_fill_2 FILLER_23_941 ();
 sg13g2_fill_1 FILLER_23_943 ();
 sg13g2_fill_1 FILLER_23_949 ();
 sg13g2_fill_1 FILLER_23_959 ();
 sg13g2_fill_1 FILLER_23_978 ();
 sg13g2_fill_1 FILLER_23_992 ();
 sg13g2_decap_4 FILLER_23_1025 ();
 sg13g2_fill_2 FILLER_24_38 ();
 sg13g2_decap_8 FILLER_24_44 ();
 sg13g2_decap_4 FILLER_24_51 ();
 sg13g2_fill_1 FILLER_24_55 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_4 FILLER_24_70 ();
 sg13g2_fill_2 FILLER_24_74 ();
 sg13g2_fill_2 FILLER_24_80 ();
 sg13g2_decap_4 FILLER_24_94 ();
 sg13g2_fill_2 FILLER_24_174 ();
 sg13g2_fill_1 FILLER_24_176 ();
 sg13g2_fill_2 FILLER_24_208 ();
 sg13g2_decap_8 FILLER_24_221 ();
 sg13g2_fill_1 FILLER_24_228 ();
 sg13g2_fill_2 FILLER_24_243 ();
 sg13g2_decap_8 FILLER_24_275 ();
 sg13g2_fill_2 FILLER_24_306 ();
 sg13g2_fill_1 FILLER_24_308 ();
 sg13g2_fill_2 FILLER_24_324 ();
 sg13g2_decap_4 FILLER_24_346 ();
 sg13g2_decap_8 FILLER_24_356 ();
 sg13g2_decap_8 FILLER_24_363 ();
 sg13g2_fill_2 FILLER_24_370 ();
 sg13g2_fill_1 FILLER_24_372 ();
 sg13g2_fill_1 FILLER_24_455 ();
 sg13g2_decap_8 FILLER_24_483 ();
 sg13g2_decap_4 FILLER_24_490 ();
 sg13g2_fill_1 FILLER_24_494 ();
 sg13g2_decap_8 FILLER_24_531 ();
 sg13g2_decap_4 FILLER_24_538 ();
 sg13g2_decap_8 FILLER_24_546 ();
 sg13g2_decap_8 FILLER_24_553 ();
 sg13g2_decap_8 FILLER_24_560 ();
 sg13g2_fill_2 FILLER_24_567 ();
 sg13g2_fill_1 FILLER_24_569 ();
 sg13g2_fill_1 FILLER_24_593 ();
 sg13g2_fill_2 FILLER_24_612 ();
 sg13g2_fill_1 FILLER_24_614 ();
 sg13g2_fill_1 FILLER_24_649 ();
 sg13g2_decap_4 FILLER_24_666 ();
 sg13g2_fill_1 FILLER_24_670 ();
 sg13g2_fill_1 FILLER_24_678 ();
 sg13g2_fill_2 FILLER_24_706 ();
 sg13g2_fill_2 FILLER_24_753 ();
 sg13g2_fill_1 FILLER_24_755 ();
 sg13g2_fill_2 FILLER_24_769 ();
 sg13g2_decap_8 FILLER_24_789 ();
 sg13g2_decap_8 FILLER_24_796 ();
 sg13g2_decap_4 FILLER_24_803 ();
 sg13g2_fill_1 FILLER_24_807 ();
 sg13g2_fill_2 FILLER_24_812 ();
 sg13g2_fill_1 FILLER_24_814 ();
 sg13g2_decap_8 FILLER_24_819 ();
 sg13g2_decap_8 FILLER_24_826 ();
 sg13g2_decap_8 FILLER_24_833 ();
 sg13g2_decap_4 FILLER_24_844 ();
 sg13g2_fill_2 FILLER_24_848 ();
 sg13g2_decap_8 FILLER_24_854 ();
 sg13g2_fill_1 FILLER_24_861 ();
 sg13g2_decap_4 FILLER_24_871 ();
 sg13g2_fill_2 FILLER_24_875 ();
 sg13g2_fill_2 FILLER_24_904 ();
 sg13g2_fill_1 FILLER_24_929 ();
 sg13g2_fill_2 FILLER_24_962 ();
 sg13g2_fill_1 FILLER_24_964 ();
 sg13g2_fill_1 FILLER_24_997 ();
 sg13g2_fill_1 FILLER_24_1007 ();
 sg13g2_decap_4 FILLER_24_1025 ();
 sg13g2_fill_1 FILLER_25_36 ();
 sg13g2_decap_8 FILLER_25_54 ();
 sg13g2_fill_2 FILLER_25_65 ();
 sg13g2_fill_1 FILLER_25_90 ();
 sg13g2_decap_4 FILLER_25_101 ();
 sg13g2_decap_8 FILLER_25_118 ();
 sg13g2_fill_1 FILLER_25_125 ();
 sg13g2_fill_2 FILLER_25_131 ();
 sg13g2_fill_2 FILLER_25_139 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_fill_1 FILLER_25_161 ();
 sg13g2_fill_2 FILLER_25_227 ();
 sg13g2_fill_2 FILLER_25_245 ();
 sg13g2_decap_8 FILLER_25_274 ();
 sg13g2_fill_2 FILLER_25_281 ();
 sg13g2_fill_1 FILLER_25_283 ();
 sg13g2_fill_2 FILLER_25_333 ();
 sg13g2_fill_1 FILLER_25_335 ();
 sg13g2_decap_8 FILLER_25_399 ();
 sg13g2_decap_8 FILLER_25_406 ();
 sg13g2_fill_1 FILLER_25_413 ();
 sg13g2_decap_4 FILLER_25_452 ();
 sg13g2_fill_2 FILLER_25_460 ();
 sg13g2_decap_8 FILLER_25_470 ();
 sg13g2_decap_8 FILLER_25_477 ();
 sg13g2_fill_1 FILLER_25_484 ();
 sg13g2_decap_8 FILLER_25_499 ();
 sg13g2_decap_8 FILLER_25_516 ();
 sg13g2_decap_8 FILLER_25_523 ();
 sg13g2_decap_4 FILLER_25_530 ();
 sg13g2_fill_2 FILLER_25_534 ();
 sg13g2_decap_8 FILLER_25_552 ();
 sg13g2_decap_8 FILLER_25_559 ();
 sg13g2_decap_4 FILLER_25_566 ();
 sg13g2_fill_2 FILLER_25_570 ();
 sg13g2_decap_8 FILLER_25_575 ();
 sg13g2_decap_8 FILLER_25_582 ();
 sg13g2_fill_1 FILLER_25_589 ();
 sg13g2_fill_2 FILLER_25_621 ();
 sg13g2_decap_8 FILLER_25_660 ();
 sg13g2_decap_8 FILLER_25_683 ();
 sg13g2_fill_2 FILLER_25_690 ();
 sg13g2_fill_1 FILLER_25_692 ();
 sg13g2_fill_2 FILLER_25_698 ();
 sg13g2_fill_1 FILLER_25_711 ();
 sg13g2_fill_2 FILLER_25_739 ();
 sg13g2_fill_1 FILLER_25_741 ();
 sg13g2_decap_4 FILLER_25_764 ();
 sg13g2_fill_2 FILLER_25_773 ();
 sg13g2_fill_1 FILLER_25_775 ();
 sg13g2_decap_4 FILLER_25_783 ();
 sg13g2_fill_2 FILLER_25_787 ();
 sg13g2_fill_1 FILLER_25_807 ();
 sg13g2_decap_8 FILLER_25_813 ();
 sg13g2_fill_1 FILLER_25_820 ();
 sg13g2_fill_2 FILLER_25_853 ();
 sg13g2_decap_4 FILLER_25_860 ();
 sg13g2_fill_2 FILLER_25_864 ();
 sg13g2_fill_2 FILLER_25_879 ();
 sg13g2_decap_4 FILLER_25_930 ();
 sg13g2_fill_2 FILLER_25_934 ();
 sg13g2_decap_4 FILLER_25_944 ();
 sg13g2_fill_2 FILLER_25_952 ();
 sg13g2_decap_8 FILLER_26_8 ();
 sg13g2_decap_8 FILLER_26_15 ();
 sg13g2_decap_4 FILLER_26_22 ();
 sg13g2_fill_1 FILLER_26_26 ();
 sg13g2_fill_1 FILLER_26_32 ();
 sg13g2_fill_2 FILLER_26_41 ();
 sg13g2_fill_1 FILLER_26_43 ();
 sg13g2_decap_4 FILLER_26_65 ();
 sg13g2_fill_1 FILLER_26_82 ();
 sg13g2_fill_2 FILLER_26_88 ();
 sg13g2_decap_8 FILLER_26_95 ();
 sg13g2_decap_4 FILLER_26_102 ();
 sg13g2_fill_1 FILLER_26_106 ();
 sg13g2_fill_2 FILLER_26_111 ();
 sg13g2_decap_8 FILLER_26_121 ();
 sg13g2_decap_8 FILLER_26_128 ();
 sg13g2_fill_2 FILLER_26_135 ();
 sg13g2_fill_1 FILLER_26_137 ();
 sg13g2_decap_8 FILLER_26_158 ();
 sg13g2_fill_1 FILLER_26_165 ();
 sg13g2_fill_2 FILLER_26_183 ();
 sg13g2_fill_1 FILLER_26_185 ();
 sg13g2_fill_2 FILLER_26_216 ();
 sg13g2_fill_1 FILLER_26_218 ();
 sg13g2_decap_8 FILLER_26_224 ();
 sg13g2_fill_2 FILLER_26_231 ();
 sg13g2_fill_2 FILLER_26_253 ();
 sg13g2_fill_1 FILLER_26_255 ();
 sg13g2_decap_8 FILLER_26_283 ();
 sg13g2_fill_1 FILLER_26_290 ();
 sg13g2_fill_2 FILLER_26_297 ();
 sg13g2_fill_1 FILLER_26_299 ();
 sg13g2_fill_1 FILLER_26_308 ();
 sg13g2_decap_8 FILLER_26_317 ();
 sg13g2_decap_8 FILLER_26_324 ();
 sg13g2_decap_8 FILLER_26_331 ();
 sg13g2_decap_4 FILLER_26_338 ();
 sg13g2_decap_4 FILLER_26_353 ();
 sg13g2_decap_8 FILLER_26_365 ();
 sg13g2_decap_8 FILLER_26_372 ();
 sg13g2_decap_8 FILLER_26_379 ();
 sg13g2_fill_1 FILLER_26_386 ();
 sg13g2_fill_1 FILLER_26_397 ();
 sg13g2_fill_2 FILLER_26_429 ();
 sg13g2_fill_2 FILLER_26_468 ();
 sg13g2_fill_1 FILLER_26_470 ();
 sg13g2_decap_8 FILLER_26_485 ();
 sg13g2_decap_8 FILLER_26_492 ();
 sg13g2_decap_4 FILLER_26_499 ();
 sg13g2_fill_1 FILLER_26_503 ();
 sg13g2_decap_8 FILLER_26_520 ();
 sg13g2_decap_4 FILLER_26_527 ();
 sg13g2_decap_8 FILLER_26_555 ();
 sg13g2_decap_4 FILLER_26_562 ();
 sg13g2_decap_4 FILLER_26_595 ();
 sg13g2_fill_1 FILLER_26_603 ();
 sg13g2_decap_8 FILLER_26_609 ();
 sg13g2_fill_1 FILLER_26_616 ();
 sg13g2_fill_1 FILLER_26_629 ();
 sg13g2_decap_4 FILLER_26_647 ();
 sg13g2_fill_2 FILLER_26_651 ();
 sg13g2_fill_2 FILLER_26_657 ();
 sg13g2_fill_1 FILLER_26_659 ();
 sg13g2_fill_2 FILLER_26_671 ();
 sg13g2_fill_1 FILLER_26_673 ();
 sg13g2_decap_8 FILLER_26_685 ();
 sg13g2_fill_2 FILLER_26_692 ();
 sg13g2_fill_1 FILLER_26_694 ();
 sg13g2_decap_4 FILLER_26_700 ();
 sg13g2_fill_1 FILLER_26_704 ();
 sg13g2_decap_8 FILLER_26_721 ();
 sg13g2_decap_4 FILLER_26_728 ();
 sg13g2_decap_8 FILLER_26_834 ();
 sg13g2_fill_1 FILLER_26_841 ();
 sg13g2_fill_1 FILLER_26_872 ();
 sg13g2_fill_1 FILLER_26_892 ();
 sg13g2_fill_2 FILLER_26_897 ();
 sg13g2_fill_1 FILLER_26_899 ();
 sg13g2_fill_1 FILLER_26_903 ();
 sg13g2_decap_8 FILLER_26_922 ();
 sg13g2_fill_2 FILLER_26_939 ();
 sg13g2_fill_1 FILLER_26_941 ();
 sg13g2_fill_2 FILLER_26_946 ();
 sg13g2_fill_1 FILLER_26_948 ();
 sg13g2_fill_2 FILLER_26_954 ();
 sg13g2_fill_2 FILLER_26_964 ();
 sg13g2_fill_1 FILLER_26_966 ();
 sg13g2_decap_8 FILLER_26_1021 ();
 sg13g2_fill_1 FILLER_26_1028 ();
 sg13g2_fill_2 FILLER_27_4 ();
 sg13g2_fill_1 FILLER_27_6 ();
 sg13g2_decap_4 FILLER_27_21 ();
 sg13g2_fill_2 FILLER_27_25 ();
 sg13g2_decap_8 FILLER_27_30 ();
 sg13g2_decap_8 FILLER_27_37 ();
 sg13g2_decap_8 FILLER_27_44 ();
 sg13g2_fill_1 FILLER_27_51 ();
 sg13g2_fill_1 FILLER_27_73 ();
 sg13g2_fill_2 FILLER_27_88 ();
 sg13g2_fill_1 FILLER_27_90 ();
 sg13g2_decap_8 FILLER_27_96 ();
 sg13g2_fill_2 FILLER_27_103 ();
 sg13g2_fill_1 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_124 ();
 sg13g2_decap_8 FILLER_27_131 ();
 sg13g2_decap_8 FILLER_27_138 ();
 sg13g2_decap_8 FILLER_27_145 ();
 sg13g2_fill_2 FILLER_27_152 ();
 sg13g2_decap_8 FILLER_27_160 ();
 sg13g2_decap_4 FILLER_27_167 ();
 sg13g2_fill_1 FILLER_27_171 ();
 sg13g2_decap_8 FILLER_27_185 ();
 sg13g2_decap_8 FILLER_27_192 ();
 sg13g2_fill_1 FILLER_27_199 ();
 sg13g2_fill_2 FILLER_27_204 ();
 sg13g2_fill_2 FILLER_27_233 ();
 sg13g2_fill_1 FILLER_27_235 ();
 sg13g2_fill_2 FILLER_27_242 ();
 sg13g2_decap_8 FILLER_27_248 ();
 sg13g2_decap_8 FILLER_27_255 ();
 sg13g2_decap_8 FILLER_27_262 ();
 sg13g2_decap_8 FILLER_27_269 ();
 sg13g2_decap_8 FILLER_27_276 ();
 sg13g2_decap_8 FILLER_27_295 ();
 sg13g2_decap_8 FILLER_27_302 ();
 sg13g2_decap_8 FILLER_27_309 ();
 sg13g2_fill_2 FILLER_27_316 ();
 sg13g2_fill_1 FILLER_27_318 ();
 sg13g2_decap_8 FILLER_27_325 ();
 sg13g2_decap_8 FILLER_27_332 ();
 sg13g2_fill_2 FILLER_27_339 ();
 sg13g2_fill_1 FILLER_27_341 ();
 sg13g2_decap_8 FILLER_27_347 ();
 sg13g2_decap_4 FILLER_27_354 ();
 sg13g2_fill_2 FILLER_27_401 ();
 sg13g2_fill_1 FILLER_27_403 ();
 sg13g2_decap_8 FILLER_27_431 ();
 sg13g2_fill_1 FILLER_27_438 ();
 sg13g2_fill_1 FILLER_27_448 ();
 sg13g2_fill_2 FILLER_27_503 ();
 sg13g2_decap_4 FILLER_27_524 ();
 sg13g2_decap_8 FILLER_27_532 ();
 sg13g2_decap_8 FILLER_27_539 ();
 sg13g2_fill_2 FILLER_27_550 ();
 sg13g2_fill_2 FILLER_27_558 ();
 sg13g2_decap_8 FILLER_27_579 ();
 sg13g2_fill_2 FILLER_27_586 ();
 sg13g2_fill_2 FILLER_27_615 ();
 sg13g2_fill_1 FILLER_27_617 ();
 sg13g2_fill_1 FILLER_27_623 ();
 sg13g2_fill_2 FILLER_27_629 ();
 sg13g2_fill_1 FILLER_27_631 ();
 sg13g2_fill_1 FILLER_27_675 ();
 sg13g2_decap_4 FILLER_27_684 ();
 sg13g2_fill_2 FILLER_27_745 ();
 sg13g2_decap_4 FILLER_27_763 ();
 sg13g2_fill_1 FILLER_27_767 ();
 sg13g2_fill_2 FILLER_27_811 ();
 sg13g2_decap_8 FILLER_27_822 ();
 sg13g2_fill_2 FILLER_27_829 ();
 sg13g2_fill_1 FILLER_27_841 ();
 sg13g2_decap_4 FILLER_27_872 ();
 sg13g2_fill_1 FILLER_27_876 ();
 sg13g2_fill_2 FILLER_27_917 ();
 sg13g2_decap_4 FILLER_27_987 ();
 sg13g2_fill_2 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_2 ();
 sg13g2_fill_1 FILLER_28_17 ();
 sg13g2_fill_2 FILLER_28_32 ();
 sg13g2_fill_2 FILLER_28_37 ();
 sg13g2_fill_1 FILLER_28_39 ();
 sg13g2_decap_4 FILLER_28_44 ();
 sg13g2_fill_1 FILLER_28_48 ();
 sg13g2_fill_2 FILLER_28_53 ();
 sg13g2_fill_1 FILLER_28_55 ();
 sg13g2_decap_4 FILLER_28_60 ();
 sg13g2_fill_2 FILLER_28_68 ();
 sg13g2_fill_1 FILLER_28_70 ();
 sg13g2_fill_2 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_94 ();
 sg13g2_decap_8 FILLER_28_101 ();
 sg13g2_fill_2 FILLER_28_108 ();
 sg13g2_fill_1 FILLER_28_110 ();
 sg13g2_decap_8 FILLER_28_132 ();
 sg13g2_decap_8 FILLER_28_150 ();
 sg13g2_decap_8 FILLER_28_157 ();
 sg13g2_decap_4 FILLER_28_164 ();
 sg13g2_decap_8 FILLER_28_177 ();
 sg13g2_decap_4 FILLER_28_184 ();
 sg13g2_fill_2 FILLER_28_188 ();
 sg13g2_decap_8 FILLER_28_199 ();
 sg13g2_decap_8 FILLER_28_206 ();
 sg13g2_decap_8 FILLER_28_213 ();
 sg13g2_decap_8 FILLER_28_220 ();
 sg13g2_fill_2 FILLER_28_227 ();
 sg13g2_decap_4 FILLER_28_251 ();
 sg13g2_fill_2 FILLER_28_261 ();
 sg13g2_fill_1 FILLER_28_263 ();
 sg13g2_decap_4 FILLER_28_273 ();
 sg13g2_fill_1 FILLER_28_277 ();
 sg13g2_fill_2 FILLER_28_292 ();
 sg13g2_decap_8 FILLER_28_302 ();
 sg13g2_fill_2 FILLER_28_332 ();
 sg13g2_fill_1 FILLER_28_334 ();
 sg13g2_decap_8 FILLER_28_355 ();
 sg13g2_fill_2 FILLER_28_362 ();
 sg13g2_decap_4 FILLER_28_374 ();
 sg13g2_decap_8 FILLER_28_382 ();
 sg13g2_decap_4 FILLER_28_408 ();
 sg13g2_fill_2 FILLER_28_446 ();
 sg13g2_fill_1 FILLER_28_448 ();
 sg13g2_decap_8 FILLER_28_470 ();
 sg13g2_decap_4 FILLER_28_477 ();
 sg13g2_fill_2 FILLER_28_485 ();
 sg13g2_fill_1 FILLER_28_487 ();
 sg13g2_decap_4 FILLER_28_493 ();
 sg13g2_fill_2 FILLER_28_497 ();
 sg13g2_fill_1 FILLER_28_503 ();
 sg13g2_fill_1 FILLER_28_509 ();
 sg13g2_decap_8 FILLER_28_547 ();
 sg13g2_decap_4 FILLER_28_554 ();
 sg13g2_fill_2 FILLER_28_566 ();
 sg13g2_fill_1 FILLER_28_568 ();
 sg13g2_fill_1 FILLER_28_592 ();
 sg13g2_decap_4 FILLER_28_597 ();
 sg13g2_fill_2 FILLER_28_601 ();
 sg13g2_decap_8 FILLER_28_612 ();
 sg13g2_fill_1 FILLER_28_619 ();
 sg13g2_decap_8 FILLER_28_634 ();
 sg13g2_fill_1 FILLER_28_641 ();
 sg13g2_decap_8 FILLER_28_659 ();
 sg13g2_fill_1 FILLER_28_666 ();
 sg13g2_fill_2 FILLER_28_687 ();
 sg13g2_fill_2 FILLER_28_748 ();
 sg13g2_fill_1 FILLER_28_769 ();
 sg13g2_fill_2 FILLER_28_777 ();
 sg13g2_fill_2 FILLER_28_783 ();
 sg13g2_fill_1 FILLER_28_785 ();
 sg13g2_fill_2 FILLER_28_789 ();
 sg13g2_fill_2 FILLER_28_800 ();
 sg13g2_fill_1 FILLER_28_806 ();
 sg13g2_decap_4 FILLER_28_834 ();
 sg13g2_fill_2 FILLER_28_871 ();
 sg13g2_decap_4 FILLER_28_877 ();
 sg13g2_fill_1 FILLER_28_881 ();
 sg13g2_decap_8 FILLER_28_886 ();
 sg13g2_decap_4 FILLER_28_893 ();
 sg13g2_fill_1 FILLER_28_902 ();
 sg13g2_fill_1 FILLER_28_946 ();
 sg13g2_decap_8 FILLER_28_960 ();
 sg13g2_decap_8 FILLER_28_967 ();
 sg13g2_decap_8 FILLER_28_974 ();
 sg13g2_decap_4 FILLER_28_981 ();
 sg13g2_fill_1 FILLER_28_985 ();
 sg13g2_fill_2 FILLER_28_1012 ();
 sg13g2_fill_1 FILLER_28_1014 ();
 sg13g2_decap_4 FILLER_28_1024 ();
 sg13g2_fill_1 FILLER_28_1028 ();
 sg13g2_decap_4 FILLER_29_4 ();
 sg13g2_decap_4 FILLER_29_17 ();
 sg13g2_fill_2 FILLER_29_27 ();
 sg13g2_decap_8 FILLER_29_32 ();
 sg13g2_decap_8 FILLER_29_65 ();
 sg13g2_decap_8 FILLER_29_72 ();
 sg13g2_decap_8 FILLER_29_79 ();
 sg13g2_fill_2 FILLER_29_86 ();
 sg13g2_fill_1 FILLER_29_88 ();
 sg13g2_fill_2 FILLER_29_104 ();
 sg13g2_fill_1 FILLER_29_106 ();
 sg13g2_decap_4 FILLER_29_111 ();
 sg13g2_fill_1 FILLER_29_115 ();
 sg13g2_fill_2 FILLER_29_129 ();
 sg13g2_fill_1 FILLER_29_131 ();
 sg13g2_fill_2 FILLER_29_167 ();
 sg13g2_fill_2 FILLER_29_258 ();
 sg13g2_fill_1 FILLER_29_260 ();
 sg13g2_decap_8 FILLER_29_269 ();
 sg13g2_fill_2 FILLER_29_276 ();
 sg13g2_fill_1 FILLER_29_278 ();
 sg13g2_decap_8 FILLER_29_302 ();
 sg13g2_decap_4 FILLER_29_309 ();
 sg13g2_decap_8 FILLER_29_318 ();
 sg13g2_decap_8 FILLER_29_325 ();
 sg13g2_decap_8 FILLER_29_332 ();
 sg13g2_fill_2 FILLER_29_339 ();
 sg13g2_decap_8 FILLER_29_351 ();
 sg13g2_decap_8 FILLER_29_358 ();
 sg13g2_decap_8 FILLER_29_365 ();
 sg13g2_decap_8 FILLER_29_372 ();
 sg13g2_decap_8 FILLER_29_379 ();
 sg13g2_fill_2 FILLER_29_386 ();
 sg13g2_decap_8 FILLER_29_415 ();
 sg13g2_decap_8 FILLER_29_422 ();
 sg13g2_decap_4 FILLER_29_471 ();
 sg13g2_decap_8 FILLER_29_507 ();
 sg13g2_fill_2 FILLER_29_514 ();
 sg13g2_decap_8 FILLER_29_563 ();
 sg13g2_decap_8 FILLER_29_570 ();
 sg13g2_fill_2 FILLER_29_577 ();
 sg13g2_fill_1 FILLER_29_605 ();
 sg13g2_fill_2 FILLER_29_710 ();
 sg13g2_fill_1 FILLER_29_717 ();
 sg13g2_fill_2 FILLER_29_797 ();
 sg13g2_fill_2 FILLER_29_848 ();
 sg13g2_fill_1 FILLER_29_858 ();
 sg13g2_fill_2 FILLER_29_895 ();
 sg13g2_fill_1 FILLER_29_897 ();
 sg13g2_fill_2 FILLER_29_960 ();
 sg13g2_fill_1 FILLER_29_962 ();
 sg13g2_fill_2 FILLER_29_969 ();
 sg13g2_decap_4 FILLER_29_977 ();
 sg13g2_fill_1 FILLER_29_981 ();
 sg13g2_fill_2 FILLER_29_1026 ();
 sg13g2_fill_1 FILLER_29_1028 ();
 sg13g2_fill_1 FILLER_30_4 ();
 sg13g2_decap_8 FILLER_30_72 ();
 sg13g2_decap_8 FILLER_30_79 ();
 sg13g2_decap_8 FILLER_30_86 ();
 sg13g2_decap_4 FILLER_30_127 ();
 sg13g2_decap_4 FILLER_30_152 ();
 sg13g2_fill_1 FILLER_30_161 ();
 sg13g2_decap_8 FILLER_30_176 ();
 sg13g2_decap_4 FILLER_30_183 ();
 sg13g2_fill_2 FILLER_30_187 ();
 sg13g2_fill_1 FILLER_30_230 ();
 sg13g2_fill_2 FILLER_30_248 ();
 sg13g2_decap_8 FILLER_30_267 ();
 sg13g2_decap_8 FILLER_30_274 ();
 sg13g2_decap_8 FILLER_30_281 ();
 sg13g2_decap_8 FILLER_30_294 ();
 sg13g2_fill_2 FILLER_30_301 ();
 sg13g2_fill_2 FILLER_30_309 ();
 sg13g2_decap_8 FILLER_30_348 ();
 sg13g2_fill_2 FILLER_30_355 ();
 sg13g2_fill_1 FILLER_30_357 ();
 sg13g2_fill_1 FILLER_30_383 ();
 sg13g2_fill_2 FILLER_30_387 ();
 sg13g2_fill_1 FILLER_30_389 ();
 sg13g2_fill_2 FILLER_30_403 ();
 sg13g2_fill_2 FILLER_30_484 ();
 sg13g2_fill_1 FILLER_30_495 ();
 sg13g2_decap_8 FILLER_30_512 ();
 sg13g2_decap_4 FILLER_30_519 ();
 sg13g2_fill_1 FILLER_30_523 ();
 sg13g2_fill_1 FILLER_30_546 ();
 sg13g2_decap_8 FILLER_30_574 ();
 sg13g2_fill_2 FILLER_30_581 ();
 sg13g2_fill_1 FILLER_30_583 ();
 sg13g2_decap_8 FILLER_30_638 ();
 sg13g2_decap_4 FILLER_30_645 ();
 sg13g2_fill_1 FILLER_30_649 ();
 sg13g2_decap_8 FILLER_30_659 ();
 sg13g2_fill_2 FILLER_30_666 ();
 sg13g2_fill_1 FILLER_30_668 ();
 sg13g2_decap_4 FILLER_30_699 ();
 sg13g2_fill_2 FILLER_30_703 ();
 sg13g2_decap_8 FILLER_30_744 ();
 sg13g2_fill_1 FILLER_30_751 ();
 sg13g2_fill_1 FILLER_30_774 ();
 sg13g2_fill_2 FILLER_30_789 ();
 sg13g2_fill_2 FILLER_30_823 ();
 sg13g2_decap_4 FILLER_30_830 ();
 sg13g2_decap_4 FILLER_30_839 ();
 sg13g2_decap_4 FILLER_30_852 ();
 sg13g2_fill_2 FILLER_30_856 ();
 sg13g2_decap_4 FILLER_30_863 ();
 sg13g2_decap_4 FILLER_30_876 ();
 sg13g2_fill_1 FILLER_30_926 ();
 sg13g2_decap_8 FILLER_30_976 ();
 sg13g2_fill_2 FILLER_30_983 ();
 sg13g2_fill_1 FILLER_30_996 ();
 sg13g2_decap_8 FILLER_31_34 ();
 sg13g2_fill_2 FILLER_31_41 ();
 sg13g2_fill_1 FILLER_31_43 ();
 sg13g2_fill_1 FILLER_31_53 ();
 sg13g2_fill_2 FILLER_31_64 ();
 sg13g2_decap_4 FILLER_31_84 ();
 sg13g2_fill_2 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_145 ();
 sg13g2_decap_8 FILLER_31_152 ();
 sg13g2_fill_1 FILLER_31_163 ();
 sg13g2_fill_2 FILLER_31_191 ();
 sg13g2_decap_4 FILLER_31_206 ();
 sg13g2_decap_8 FILLER_31_213 ();
 sg13g2_decap_8 FILLER_31_220 ();
 sg13g2_decap_8 FILLER_31_227 ();
 sg13g2_decap_8 FILLER_31_234 ();
 sg13g2_decap_8 FILLER_31_241 ();
 sg13g2_decap_8 FILLER_31_248 ();
 sg13g2_fill_2 FILLER_31_255 ();
 sg13g2_fill_1 FILLER_31_257 ();
 sg13g2_decap_8 FILLER_31_264 ();
 sg13g2_decap_8 FILLER_31_271 ();
 sg13g2_decap_4 FILLER_31_278 ();
 sg13g2_fill_2 FILLER_31_282 ();
 sg13g2_decap_8 FILLER_31_288 ();
 sg13g2_decap_8 FILLER_31_295 ();
 sg13g2_decap_8 FILLER_31_302 ();
 sg13g2_decap_4 FILLER_31_309 ();
 sg13g2_decap_8 FILLER_31_317 ();
 sg13g2_fill_1 FILLER_31_324 ();
 sg13g2_decap_8 FILLER_31_331 ();
 sg13g2_decap_8 FILLER_31_338 ();
 sg13g2_decap_4 FILLER_31_345 ();
 sg13g2_fill_1 FILLER_31_349 ();
 sg13g2_decap_4 FILLER_31_355 ();
 sg13g2_fill_1 FILLER_31_359 ();
 sg13g2_decap_4 FILLER_31_387 ();
 sg13g2_fill_2 FILLER_31_391 ();
 sg13g2_decap_8 FILLER_31_403 ();
 sg13g2_fill_2 FILLER_31_410 ();
 sg13g2_fill_1 FILLER_31_412 ();
 sg13g2_fill_2 FILLER_31_468 ();
 sg13g2_fill_1 FILLER_31_470 ();
 sg13g2_decap_4 FILLER_31_480 ();
 sg13g2_decap_8 FILLER_31_501 ();
 sg13g2_decap_4 FILLER_31_508 ();
 sg13g2_fill_1 FILLER_31_512 ();
 sg13g2_decap_4 FILLER_31_516 ();
 sg13g2_fill_1 FILLER_31_525 ();
 sg13g2_decap_8 FILLER_31_538 ();
 sg13g2_decap_8 FILLER_31_545 ();
 sg13g2_decap_8 FILLER_31_552 ();
 sg13g2_fill_1 FILLER_31_559 ();
 sg13g2_decap_8 FILLER_31_591 ();
 sg13g2_decap_4 FILLER_31_606 ();
 sg13g2_fill_1 FILLER_31_610 ();
 sg13g2_decap_4 FILLER_31_619 ();
 sg13g2_fill_2 FILLER_31_623 ();
 sg13g2_fill_2 FILLER_31_638 ();
 sg13g2_fill_2 FILLER_31_645 ();
 sg13g2_decap_8 FILLER_31_652 ();
 sg13g2_fill_2 FILLER_31_659 ();
 sg13g2_fill_2 FILLER_31_669 ();
 sg13g2_fill_1 FILLER_31_671 ();
 sg13g2_fill_1 FILLER_31_690 ();
 sg13g2_fill_1 FILLER_31_696 ();
 sg13g2_fill_1 FILLER_31_710 ();
 sg13g2_fill_2 FILLER_31_724 ();
 sg13g2_fill_1 FILLER_31_726 ();
 sg13g2_fill_2 FILLER_31_732 ();
 sg13g2_fill_1 FILLER_31_734 ();
 sg13g2_decap_8 FILLER_31_740 ();
 sg13g2_decap_4 FILLER_31_747 ();
 sg13g2_fill_2 FILLER_31_805 ();
 sg13g2_fill_1 FILLER_31_816 ();
 sg13g2_fill_2 FILLER_31_823 ();
 sg13g2_decap_4 FILLER_31_834 ();
 sg13g2_fill_1 FILLER_31_838 ();
 sg13g2_fill_1 FILLER_31_861 ();
 sg13g2_fill_2 FILLER_31_921 ();
 sg13g2_fill_1 FILLER_31_965 ();
 sg13g2_decap_8 FILLER_32_31 ();
 sg13g2_decap_4 FILLER_32_38 ();
 sg13g2_fill_1 FILLER_32_42 ();
 sg13g2_decap_4 FILLER_32_72 ();
 sg13g2_fill_1 FILLER_32_76 ();
 sg13g2_decap_8 FILLER_32_121 ();
 sg13g2_fill_2 FILLER_32_128 ();
 sg13g2_fill_2 FILLER_32_144 ();
 sg13g2_fill_1 FILLER_32_146 ();
 sg13g2_fill_2 FILLER_32_173 ();
 sg13g2_fill_1 FILLER_32_205 ();
 sg13g2_decap_8 FILLER_32_211 ();
 sg13g2_decap_8 FILLER_32_218 ();
 sg13g2_fill_1 FILLER_32_233 ();
 sg13g2_decap_8 FILLER_32_240 ();
 sg13g2_decap_4 FILLER_32_247 ();
 sg13g2_fill_1 FILLER_32_251 ();
 sg13g2_fill_1 FILLER_32_263 ();
 sg13g2_decap_8 FILLER_32_269 ();
 sg13g2_decap_4 FILLER_32_276 ();
 sg13g2_decap_4 FILLER_32_296 ();
 sg13g2_decap_8 FILLER_32_306 ();
 sg13g2_decap_8 FILLER_32_313 ();
 sg13g2_fill_2 FILLER_32_320 ();
 sg13g2_decap_4 FILLER_32_338 ();
 sg13g2_decap_8 FILLER_32_357 ();
 sg13g2_fill_2 FILLER_32_364 ();
 sg13g2_fill_2 FILLER_32_391 ();
 sg13g2_fill_1 FILLER_32_393 ();
 sg13g2_fill_1 FILLER_32_404 ();
 sg13g2_fill_1 FILLER_32_432 ();
 sg13g2_fill_2 FILLER_32_460 ();
 sg13g2_decap_4 FILLER_32_498 ();
 sg13g2_fill_2 FILLER_32_566 ();
 sg13g2_fill_2 FILLER_32_577 ();
 sg13g2_fill_2 FILLER_32_606 ();
 sg13g2_decap_4 FILLER_32_628 ();
 sg13g2_fill_2 FILLER_32_632 ();
 sg13g2_decap_8 FILLER_32_755 ();
 sg13g2_fill_2 FILLER_32_762 ();
 sg13g2_fill_2 FILLER_32_818 ();
 sg13g2_fill_1 FILLER_32_820 ();
 sg13g2_fill_2 FILLER_32_826 ();
 sg13g2_fill_2 FILLER_32_833 ();
 sg13g2_fill_1 FILLER_32_835 ();
 sg13g2_decap_8 FILLER_32_853 ();
 sg13g2_fill_1 FILLER_32_860 ();
 sg13g2_fill_1 FILLER_32_901 ();
 sg13g2_fill_2 FILLER_32_907 ();
 sg13g2_fill_2 FILLER_32_918 ();
 sg13g2_fill_1 FILLER_32_920 ();
 sg13g2_fill_2 FILLER_32_975 ();
 sg13g2_fill_2 FILLER_32_983 ();
 sg13g2_decap_8 FILLER_33_4 ();
 sg13g2_fill_2 FILLER_33_11 ();
 sg13g2_fill_1 FILLER_33_23 ();
 sg13g2_fill_2 FILLER_33_54 ();
 sg13g2_fill_1 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_69 ();
 sg13g2_decap_4 FILLER_33_76 ();
 sg13g2_fill_2 FILLER_33_80 ();
 sg13g2_fill_2 FILLER_33_114 ();
 sg13g2_decap_8 FILLER_33_121 ();
 sg13g2_decap_8 FILLER_33_128 ();
 sg13g2_decap_8 FILLER_33_139 ();
 sg13g2_decap_8 FILLER_33_146 ();
 sg13g2_decap_8 FILLER_33_153 ();
 sg13g2_fill_2 FILLER_33_160 ();
 sg13g2_fill_1 FILLER_33_162 ();
 sg13g2_fill_2 FILLER_33_247 ();
 sg13g2_fill_2 FILLER_33_273 ();
 sg13g2_fill_1 FILLER_33_275 ();
 sg13g2_fill_2 FILLER_33_306 ();
 sg13g2_fill_1 FILLER_33_308 ();
 sg13g2_fill_2 FILLER_33_325 ();
 sg13g2_fill_1 FILLER_33_327 ();
 sg13g2_fill_1 FILLER_33_334 ();
 sg13g2_fill_2 FILLER_33_361 ();
 sg13g2_decap_4 FILLER_33_400 ();
 sg13g2_fill_1 FILLER_33_431 ();
 sg13g2_decap_8 FILLER_33_506 ();
 sg13g2_decap_4 FILLER_33_513 ();
 sg13g2_fill_2 FILLER_33_517 ();
 sg13g2_fill_2 FILLER_33_528 ();
 sg13g2_decap_8 FILLER_33_548 ();
 sg13g2_decap_4 FILLER_33_555 ();
 sg13g2_fill_1 FILLER_33_559 ();
 sg13g2_decap_4 FILLER_33_575 ();
 sg13g2_fill_1 FILLER_33_579 ();
 sg13g2_fill_2 FILLER_33_589 ();
 sg13g2_fill_1 FILLER_33_591 ();
 sg13g2_decap_4 FILLER_33_629 ();
 sg13g2_fill_1 FILLER_33_633 ();
 sg13g2_decap_8 FILLER_33_643 ();
 sg13g2_fill_2 FILLER_33_650 ();
 sg13g2_fill_1 FILLER_33_652 ();
 sg13g2_fill_1 FILLER_33_680 ();
 sg13g2_fill_2 FILLER_33_688 ();
 sg13g2_fill_1 FILLER_33_690 ();
 sg13g2_decap_4 FILLER_33_705 ();
 sg13g2_decap_8 FILLER_33_744 ();
 sg13g2_decap_4 FILLER_33_751 ();
 sg13g2_fill_1 FILLER_33_755 ();
 sg13g2_decap_8 FILLER_33_761 ();
 sg13g2_fill_1 FILLER_33_780 ();
 sg13g2_decap_4 FILLER_33_786 ();
 sg13g2_fill_2 FILLER_33_790 ();
 sg13g2_decap_8 FILLER_33_805 ();
 sg13g2_fill_1 FILLER_33_830 ();
 sg13g2_fill_2 FILLER_33_838 ();
 sg13g2_decap_8 FILLER_33_850 ();
 sg13g2_fill_2 FILLER_33_857 ();
 sg13g2_fill_1 FILLER_33_859 ();
 sg13g2_fill_2 FILLER_33_904 ();
 sg13g2_fill_1 FILLER_33_906 ();
 sg13g2_fill_1 FILLER_33_949 ();
 sg13g2_fill_1 FILLER_33_978 ();
 sg13g2_fill_1 FILLER_33_988 ();
 sg13g2_fill_1 FILLER_33_994 ();
 sg13g2_fill_2 FILLER_33_1027 ();
 sg13g2_fill_2 FILLER_34_4 ();
 sg13g2_fill_1 FILLER_34_6 ();
 sg13g2_decap_8 FILLER_34_29 ();
 sg13g2_decap_8 FILLER_34_36 ();
 sg13g2_decap_8 FILLER_34_43 ();
 sg13g2_decap_4 FILLER_34_50 ();
 sg13g2_decap_8 FILLER_34_80 ();
 sg13g2_decap_8 FILLER_34_87 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_4 FILLER_34_110 ();
 sg13g2_decap_4 FILLER_34_124 ();
 sg13g2_decap_4 FILLER_34_133 ();
 sg13g2_fill_1 FILLER_34_137 ();
 sg13g2_fill_2 FILLER_34_145 ();
 sg13g2_fill_1 FILLER_34_147 ();
 sg13g2_fill_1 FILLER_34_152 ();
 sg13g2_decap_4 FILLER_34_157 ();
 sg13g2_fill_2 FILLER_34_161 ();
 sg13g2_fill_2 FILLER_34_168 ();
 sg13g2_fill_1 FILLER_34_170 ();
 sg13g2_decap_8 FILLER_34_174 ();
 sg13g2_decap_4 FILLER_34_181 ();
 sg13g2_fill_1 FILLER_34_185 ();
 sg13g2_fill_2 FILLER_34_208 ();
 sg13g2_decap_8 FILLER_34_214 ();
 sg13g2_fill_2 FILLER_34_221 ();
 sg13g2_decap_8 FILLER_34_241 ();
 sg13g2_decap_8 FILLER_34_248 ();
 sg13g2_fill_2 FILLER_34_255 ();
 sg13g2_fill_1 FILLER_34_257 ();
 sg13g2_decap_8 FILLER_34_264 ();
 sg13g2_decap_8 FILLER_34_271 ();
 sg13g2_fill_2 FILLER_34_278 ();
 sg13g2_decap_8 FILLER_34_293 ();
 sg13g2_fill_2 FILLER_34_300 ();
 sg13g2_fill_1 FILLER_34_302 ();
 sg13g2_decap_8 FILLER_34_308 ();
 sg13g2_decap_4 FILLER_34_315 ();
 sg13g2_decap_8 FILLER_34_331 ();
 sg13g2_decap_8 FILLER_34_338 ();
 sg13g2_fill_2 FILLER_34_353 ();
 sg13g2_fill_1 FILLER_34_359 ();
 sg13g2_fill_1 FILLER_34_397 ();
 sg13g2_fill_2 FILLER_34_433 ();
 sg13g2_fill_1 FILLER_34_471 ();
 sg13g2_decap_8 FILLER_34_507 ();
 sg13g2_decap_8 FILLER_34_514 ();
 sg13g2_decap_8 FILLER_34_542 ();
 sg13g2_decap_4 FILLER_34_549 ();
 sg13g2_fill_2 FILLER_34_553 ();
 sg13g2_decap_4 FILLER_34_623 ();
 sg13g2_fill_1 FILLER_34_627 ();
 sg13g2_fill_2 FILLER_34_669 ();
 sg13g2_fill_1 FILLER_34_671 ();
 sg13g2_fill_1 FILLER_34_677 ();
 sg13g2_decap_8 FILLER_34_714 ();
 sg13g2_fill_2 FILLER_34_736 ();
 sg13g2_fill_1 FILLER_34_765 ();
 sg13g2_fill_1 FILLER_34_795 ();
 sg13g2_fill_2 FILLER_34_800 ();
 sg13g2_fill_1 FILLER_34_811 ();
 sg13g2_decap_8 FILLER_34_825 ();
 sg13g2_decap_8 FILLER_34_832 ();
 sg13g2_decap_4 FILLER_34_839 ();
 sg13g2_fill_2 FILLER_34_843 ();
 sg13g2_decap_4 FILLER_34_849 ();
 sg13g2_fill_1 FILLER_34_853 ();
 sg13g2_fill_2 FILLER_34_859 ();
 sg13g2_fill_2 FILLER_34_929 ();
 sg13g2_fill_1 FILLER_34_931 ();
 sg13g2_fill_1 FILLER_34_989 ();
 sg13g2_decap_4 FILLER_35_4 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_fill_2 FILLER_35_42 ();
 sg13g2_fill_1 FILLER_35_59 ();
 sg13g2_fill_2 FILLER_35_73 ();
 sg13g2_fill_2 FILLER_35_80 ();
 sg13g2_fill_1 FILLER_35_82 ();
 sg13g2_fill_1 FILLER_35_101 ();
 sg13g2_decap_4 FILLER_35_108 ();
 sg13g2_fill_2 FILLER_35_112 ();
 sg13g2_fill_1 FILLER_35_194 ();
 sg13g2_fill_2 FILLER_35_200 ();
 sg13g2_decap_8 FILLER_35_229 ();
 sg13g2_fill_1 FILLER_35_236 ();
 sg13g2_fill_2 FILLER_35_242 ();
 sg13g2_fill_1 FILLER_35_244 ();
 sg13g2_fill_2 FILLER_35_249 ();
 sg13g2_fill_1 FILLER_35_251 ();
 sg13g2_fill_1 FILLER_35_258 ();
 sg13g2_fill_1 FILLER_35_265 ();
 sg13g2_decap_8 FILLER_35_271 ();
 sg13g2_decap_8 FILLER_35_278 ();
 sg13g2_decap_8 FILLER_35_295 ();
 sg13g2_decap_8 FILLER_35_314 ();
 sg13g2_fill_2 FILLER_35_321 ();
 sg13g2_decap_8 FILLER_35_327 ();
 sg13g2_decap_8 FILLER_35_334 ();
 sg13g2_decap_4 FILLER_35_341 ();
 sg13g2_decap_4 FILLER_35_352 ();
 sg13g2_decap_4 FILLER_35_363 ();
 sg13g2_fill_1 FILLER_35_367 ();
 sg13g2_decap_8 FILLER_35_372 ();
 sg13g2_decap_8 FILLER_35_379 ();
 sg13g2_decap_8 FILLER_35_386 ();
 sg13g2_fill_2 FILLER_35_393 ();
 sg13g2_fill_1 FILLER_35_418 ();
 sg13g2_fill_2 FILLER_35_435 ();
 sg13g2_fill_1 FILLER_35_458 ();
 sg13g2_fill_2 FILLER_35_486 ();
 sg13g2_fill_1 FILLER_35_488 ();
 sg13g2_fill_1 FILLER_35_505 ();
 sg13g2_fill_2 FILLER_35_511 ();
 sg13g2_fill_1 FILLER_35_513 ();
 sg13g2_decap_4 FILLER_35_524 ();
 sg13g2_fill_1 FILLER_35_528 ();
 sg13g2_decap_8 FILLER_35_538 ();
 sg13g2_decap_8 FILLER_35_545 ();
 sg13g2_decap_4 FILLER_35_573 ();
 sg13g2_fill_2 FILLER_35_577 ();
 sg13g2_decap_4 FILLER_35_596 ();
 sg13g2_fill_2 FILLER_35_658 ();
 sg13g2_fill_1 FILLER_35_692 ();
 sg13g2_decap_8 FILLER_35_707 ();
 sg13g2_fill_2 FILLER_35_714 ();
 sg13g2_decap_4 FILLER_35_723 ();
 sg13g2_fill_2 FILLER_35_727 ();
 sg13g2_decap_8 FILLER_35_816 ();
 sg13g2_fill_2 FILLER_35_832 ();
 sg13g2_fill_1 FILLER_35_834 ();
 sg13g2_fill_1 FILLER_35_867 ();
 sg13g2_decap_4 FILLER_35_887 ();
 sg13g2_fill_1 FILLER_35_891 ();
 sg13g2_fill_1 FILLER_35_904 ();
 sg13g2_fill_1 FILLER_35_914 ();
 sg13g2_fill_2 FILLER_35_941 ();
 sg13g2_fill_2 FILLER_36_4 ();
 sg13g2_fill_1 FILLER_36_6 ();
 sg13g2_fill_2 FILLER_36_17 ();
 sg13g2_fill_1 FILLER_36_19 ();
 sg13g2_fill_1 FILLER_36_55 ();
 sg13g2_decap_4 FILLER_36_63 ();
 sg13g2_fill_2 FILLER_36_67 ();
 sg13g2_fill_2 FILLER_36_76 ();
 sg13g2_fill_2 FILLER_36_99 ();
 sg13g2_fill_1 FILLER_36_101 ();
 sg13g2_decap_4 FILLER_36_134 ();
 sg13g2_fill_2 FILLER_36_138 ();
 sg13g2_decap_4 FILLER_36_155 ();
 sg13g2_fill_1 FILLER_36_159 ();
 sg13g2_fill_2 FILLER_36_169 ();
 sg13g2_fill_1 FILLER_36_171 ();
 sg13g2_fill_1 FILLER_36_176 ();
 sg13g2_fill_2 FILLER_36_192 ();
 sg13g2_fill_1 FILLER_36_230 ();
 sg13g2_decap_4 FILLER_36_272 ();
 sg13g2_fill_2 FILLER_36_276 ();
 sg13g2_fill_2 FILLER_36_297 ();
 sg13g2_fill_1 FILLER_36_299 ();
 sg13g2_fill_2 FILLER_36_332 ();
 sg13g2_fill_1 FILLER_36_334 ();
 sg13g2_decap_8 FILLER_36_371 ();
 sg13g2_decap_8 FILLER_36_378 ();
 sg13g2_fill_1 FILLER_36_385 ();
 sg13g2_fill_2 FILLER_36_423 ();
 sg13g2_fill_2 FILLER_36_457 ();
 sg13g2_fill_1 FILLER_36_459 ();
 sg13g2_fill_2 FILLER_36_487 ();
 sg13g2_fill_1 FILLER_36_489 ();
 sg13g2_fill_2 FILLER_36_517 ();
 sg13g2_decap_4 FILLER_36_550 ();
 sg13g2_fill_1 FILLER_36_554 ();
 sg13g2_decap_8 FILLER_36_560 ();
 sg13g2_fill_2 FILLER_36_567 ();
 sg13g2_fill_2 FILLER_36_579 ();
 sg13g2_fill_1 FILLER_36_581 ();
 sg13g2_decap_8 FILLER_36_599 ();
 sg13g2_fill_1 FILLER_36_606 ();
 sg13g2_fill_2 FILLER_36_624 ();
 sg13g2_fill_1 FILLER_36_626 ();
 sg13g2_fill_1 FILLER_36_647 ();
 sg13g2_decap_4 FILLER_36_678 ();
 sg13g2_fill_1 FILLER_36_717 ();
 sg13g2_decap_8 FILLER_36_732 ();
 sg13g2_fill_2 FILLER_36_761 ();
 sg13g2_fill_2 FILLER_36_773 ();
 sg13g2_fill_2 FILLER_36_791 ();
 sg13g2_fill_1 FILLER_36_793 ();
 sg13g2_fill_2 FILLER_36_825 ();
 sg13g2_fill_1 FILLER_36_827 ();
 sg13g2_fill_1 FILLER_36_833 ();
 sg13g2_decap_4 FILLER_36_852 ();
 sg13g2_fill_1 FILLER_36_856 ();
 sg13g2_fill_1 FILLER_36_874 ();
 sg13g2_fill_2 FILLER_36_886 ();
 sg13g2_fill_2 FILLER_36_933 ();
 sg13g2_fill_1 FILLER_36_994 ();
 sg13g2_fill_1 FILLER_36_1000 ();
 sg13g2_fill_1 FILLER_36_1028 ();
 sg13g2_fill_2 FILLER_37_4 ();
 sg13g2_fill_1 FILLER_37_6 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_fill_2 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_37 ();
 sg13g2_decap_4 FILLER_37_44 ();
 sg13g2_fill_1 FILLER_37_48 ();
 sg13g2_decap_4 FILLER_37_55 ();
 sg13g2_decap_8 FILLER_37_64 ();
 sg13g2_decap_8 FILLER_37_71 ();
 sg13g2_fill_1 FILLER_37_78 ();
 sg13g2_fill_1 FILLER_37_83 ();
 sg13g2_decap_4 FILLER_37_90 ();
 sg13g2_fill_1 FILLER_37_94 ();
 sg13g2_fill_2 FILLER_37_103 ();
 sg13g2_decap_8 FILLER_37_114 ();
 sg13g2_decap_4 FILLER_37_121 ();
 sg13g2_fill_2 FILLER_37_125 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_4 FILLER_37_147 ();
 sg13g2_decap_4 FILLER_37_169 ();
 sg13g2_fill_1 FILLER_37_173 ();
 sg13g2_decap_8 FILLER_37_240 ();
 sg13g2_decap_8 FILLER_37_247 ();
 sg13g2_decap_8 FILLER_37_254 ();
 sg13g2_decap_8 FILLER_37_264 ();
 sg13g2_decap_8 FILLER_37_271 ();
 sg13g2_decap_4 FILLER_37_278 ();
 sg13g2_fill_2 FILLER_37_282 ();
 sg13g2_fill_2 FILLER_37_298 ();
 sg13g2_fill_2 FILLER_37_312 ();
 sg13g2_fill_1 FILLER_37_314 ();
 sg13g2_decap_8 FILLER_37_323 ();
 sg13g2_fill_2 FILLER_37_330 ();
 sg13g2_fill_1 FILLER_37_332 ();
 sg13g2_decap_8 FILLER_37_356 ();
 sg13g2_decap_8 FILLER_37_363 ();
 sg13g2_fill_2 FILLER_37_370 ();
 sg13g2_fill_1 FILLER_37_372 ();
 sg13g2_fill_2 FILLER_37_467 ();
 sg13g2_fill_1 FILLER_37_496 ();
 sg13g2_fill_1 FILLER_37_502 ();
 sg13g2_fill_1 FILLER_37_517 ();
 sg13g2_decap_8 FILLER_37_541 ();
 sg13g2_decap_8 FILLER_37_564 ();
 sg13g2_fill_2 FILLER_37_571 ();
 sg13g2_fill_2 FILLER_37_578 ();
 sg13g2_decap_4 FILLER_37_587 ();
 sg13g2_decap_8 FILLER_37_618 ();
 sg13g2_decap_4 FILLER_37_625 ();
 sg13g2_fill_1 FILLER_37_629 ();
 sg13g2_decap_8 FILLER_37_679 ();
 sg13g2_decap_8 FILLER_37_686 ();
 sg13g2_fill_2 FILLER_37_711 ();
 sg13g2_fill_1 FILLER_37_781 ();
 sg13g2_fill_2 FILLER_37_796 ();
 sg13g2_fill_2 FILLER_37_819 ();
 sg13g2_decap_4 FILLER_37_901 ();
 sg13g2_fill_2 FILLER_37_954 ();
 sg13g2_fill_1 FILLER_37_960 ();
 sg13g2_fill_2 FILLER_37_970 ();
 sg13g2_fill_1 FILLER_37_972 ();
 sg13g2_fill_1 FILLER_37_982 ();
 sg13g2_fill_1 FILLER_37_1001 ();
 sg13g2_fill_2 FILLER_37_1011 ();
 sg13g2_fill_2 FILLER_37_1026 ();
 sg13g2_fill_1 FILLER_37_1028 ();
 sg13g2_fill_2 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_2 ();
 sg13g2_decap_4 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_fill_2 FILLER_38_63 ();
 sg13g2_fill_1 FILLER_38_65 ();
 sg13g2_decap_8 FILLER_38_93 ();
 sg13g2_fill_2 FILLER_38_100 ();
 sg13g2_fill_1 FILLER_38_102 ();
 sg13g2_decap_8 FILLER_38_118 ();
 sg13g2_decap_8 FILLER_38_125 ();
 sg13g2_fill_2 FILLER_38_132 ();
 sg13g2_fill_1 FILLER_38_143 ();
 sg13g2_decap_8 FILLER_38_154 ();
 sg13g2_fill_2 FILLER_38_161 ();
 sg13g2_fill_1 FILLER_38_163 ();
 sg13g2_decap_8 FILLER_38_172 ();
 sg13g2_fill_2 FILLER_38_179 ();
 sg13g2_fill_1 FILLER_38_181 ();
 sg13g2_fill_1 FILLER_38_188 ();
 sg13g2_decap_4 FILLER_38_193 ();
 sg13g2_fill_1 FILLER_38_202 ();
 sg13g2_decap_8 FILLER_38_241 ();
 sg13g2_fill_1 FILLER_38_248 ();
 sg13g2_decap_4 FILLER_38_281 ();
 sg13g2_fill_2 FILLER_38_285 ();
 sg13g2_decap_8 FILLER_38_293 ();
 sg13g2_fill_2 FILLER_38_300 ();
 sg13g2_fill_1 FILLER_38_302 ();
 sg13g2_fill_1 FILLER_38_309 ();
 sg13g2_decap_8 FILLER_38_315 ();
 sg13g2_decap_8 FILLER_38_322 ();
 sg13g2_decap_8 FILLER_38_329 ();
 sg13g2_decap_4 FILLER_38_336 ();
 sg13g2_fill_2 FILLER_38_340 ();
 sg13g2_decap_4 FILLER_38_347 ();
 sg13g2_fill_1 FILLER_38_357 ();
 sg13g2_fill_2 FILLER_38_401 ();
 sg13g2_fill_2 FILLER_38_430 ();
 sg13g2_fill_2 FILLER_38_490 ();
 sg13g2_fill_1 FILLER_38_492 ();
 sg13g2_fill_1 FILLER_38_511 ();
 sg13g2_fill_1 FILLER_38_521 ();
 sg13g2_fill_1 FILLER_38_549 ();
 sg13g2_decap_8 FILLER_38_570 ();
 sg13g2_decap_8 FILLER_38_577 ();
 sg13g2_fill_1 FILLER_38_584 ();
 sg13g2_fill_2 FILLER_38_590 ();
 sg13g2_decap_4 FILLER_38_610 ();
 sg13g2_fill_1 FILLER_38_688 ();
 sg13g2_fill_1 FILLER_38_698 ();
 sg13g2_fill_2 FILLER_38_707 ();
 sg13g2_fill_1 FILLER_38_709 ();
 sg13g2_fill_1 FILLER_38_717 ();
 sg13g2_decap_8 FILLER_38_736 ();
 sg13g2_decap_4 FILLER_38_743 ();
 sg13g2_fill_1 FILLER_38_751 ();
 sg13g2_fill_1 FILLER_38_793 ();
 sg13g2_fill_1 FILLER_38_798 ();
 sg13g2_fill_2 FILLER_38_835 ();
 sg13g2_fill_2 FILLER_38_864 ();
 sg13g2_fill_1 FILLER_38_880 ();
 sg13g2_decap_8 FILLER_38_891 ();
 sg13g2_decap_8 FILLER_38_898 ();
 sg13g2_decap_8 FILLER_38_905 ();
 sg13g2_fill_2 FILLER_38_912 ();
 sg13g2_fill_1 FILLER_38_927 ();
 sg13g2_fill_2 FILLER_38_957 ();
 sg13g2_fill_1 FILLER_38_959 ();
 sg13g2_fill_1 FILLER_38_996 ();
 sg13g2_fill_1 FILLER_39_0 ();
 sg13g2_fill_2 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_57 ();
 sg13g2_fill_2 FILLER_39_75 ();
 sg13g2_fill_1 FILLER_39_85 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_decap_4 FILLER_39_98 ();
 sg13g2_fill_2 FILLER_39_102 ();
 sg13g2_decap_8 FILLER_39_109 ();
 sg13g2_decap_8 FILLER_39_116 ();
 sg13g2_fill_2 FILLER_39_123 ();
 sg13g2_fill_2 FILLER_39_135 ();
 sg13g2_fill_1 FILLER_39_150 ();
 sg13g2_decap_8 FILLER_39_157 ();
 sg13g2_fill_1 FILLER_39_164 ();
 sg13g2_decap_4 FILLER_39_170 ();
 sg13g2_decap_8 FILLER_39_179 ();
 sg13g2_fill_2 FILLER_39_186 ();
 sg13g2_fill_2 FILLER_39_195 ();
 sg13g2_decap_8 FILLER_39_205 ();
 sg13g2_fill_2 FILLER_39_212 ();
 sg13g2_fill_1 FILLER_39_214 ();
 sg13g2_decap_8 FILLER_39_239 ();
 sg13g2_decap_8 FILLER_39_246 ();
 sg13g2_decap_8 FILLER_39_253 ();
 sg13g2_decap_8 FILLER_39_260 ();
 sg13g2_decap_8 FILLER_39_267 ();
 sg13g2_decap_4 FILLER_39_274 ();
 sg13g2_fill_1 FILLER_39_278 ();
 sg13g2_fill_1 FILLER_39_284 ();
 sg13g2_decap_8 FILLER_39_302 ();
 sg13g2_decap_4 FILLER_39_309 ();
 sg13g2_fill_2 FILLER_39_313 ();
 sg13g2_decap_4 FILLER_39_321 ();
 sg13g2_decap_8 FILLER_39_337 ();
 sg13g2_fill_1 FILLER_39_344 ();
 sg13g2_fill_2 FILLER_39_360 ();
 sg13g2_decap_8 FILLER_39_366 ();
 sg13g2_decap_8 FILLER_39_373 ();
 sg13g2_decap_8 FILLER_39_423 ();
 sg13g2_decap_4 FILLER_39_430 ();
 sg13g2_fill_1 FILLER_39_434 ();
 sg13g2_fill_2 FILLER_39_465 ();
 sg13g2_fill_1 FILLER_39_516 ();
 sg13g2_decap_4 FILLER_39_535 ();
 sg13g2_fill_1 FILLER_39_560 ();
 sg13g2_decap_4 FILLER_39_588 ();
 sg13g2_fill_1 FILLER_39_592 ();
 sg13g2_fill_2 FILLER_39_654 ();
 sg13g2_fill_2 FILLER_39_664 ();
 sg13g2_decap_4 FILLER_39_705 ();
 sg13g2_fill_2 FILLER_39_709 ();
 sg13g2_fill_2 FILLER_39_725 ();
 sg13g2_fill_2 FILLER_39_779 ();
 sg13g2_fill_1 FILLER_39_790 ();
 sg13g2_fill_1 FILLER_39_858 ();
 sg13g2_fill_1 FILLER_39_864 ();
 sg13g2_fill_1 FILLER_39_878 ();
 sg13g2_fill_2 FILLER_39_911 ();
 sg13g2_fill_1 FILLER_39_913 ();
 sg13g2_fill_2 FILLER_39_969 ();
 sg13g2_fill_1 FILLER_39_971 ();
 sg13g2_fill_1 FILLER_39_977 ();
 sg13g2_fill_2 FILLER_39_983 ();
 sg13g2_fill_1 FILLER_39_985 ();
 sg13g2_fill_2 FILLER_39_1015 ();
 sg13g2_fill_1 FILLER_39_1017 ();
 sg13g2_fill_2 FILLER_39_1027 ();
 sg13g2_decap_4 FILLER_40_8 ();
 sg13g2_fill_1 FILLER_40_29 ();
 sg13g2_fill_2 FILLER_40_36 ();
 sg13g2_fill_1 FILLER_40_38 ();
 sg13g2_fill_1 FILLER_40_48 ();
 sg13g2_decap_4 FILLER_40_82 ();
 sg13g2_decap_4 FILLER_40_94 ();
 sg13g2_fill_2 FILLER_40_98 ();
 sg13g2_decap_8 FILLER_40_120 ();
 sg13g2_fill_2 FILLER_40_127 ();
 sg13g2_fill_1 FILLER_40_129 ();
 sg13g2_decap_8 FILLER_40_135 ();
 sg13g2_fill_1 FILLER_40_142 ();
 sg13g2_fill_2 FILLER_40_162 ();
 sg13g2_fill_1 FILLER_40_164 ();
 sg13g2_decap_8 FILLER_40_175 ();
 sg13g2_fill_1 FILLER_40_219 ();
 sg13g2_decap_8 FILLER_40_231 ();
 sg13g2_decap_8 FILLER_40_238 ();
 sg13g2_fill_1 FILLER_40_245 ();
 sg13g2_decap_8 FILLER_40_265 ();
 sg13g2_decap_4 FILLER_40_272 ();
 sg13g2_fill_2 FILLER_40_276 ();
 sg13g2_decap_8 FILLER_40_300 ();
 sg13g2_fill_2 FILLER_40_307 ();
 sg13g2_fill_1 FILLER_40_309 ();
 sg13g2_fill_2 FILLER_40_322 ();
 sg13g2_decap_8 FILLER_40_336 ();
 sg13g2_decap_8 FILLER_40_343 ();
 sg13g2_decap_4 FILLER_40_350 ();
 sg13g2_fill_1 FILLER_40_354 ();
 sg13g2_decap_8 FILLER_40_365 ();
 sg13g2_fill_1 FILLER_40_372 ();
 sg13g2_decap_4 FILLER_40_393 ();
 sg13g2_fill_1 FILLER_40_455 ();
 sg13g2_fill_2 FILLER_40_460 ();
 sg13g2_fill_1 FILLER_40_462 ();
 sg13g2_fill_2 FILLER_40_471 ();
 sg13g2_decap_8 FILLER_40_477 ();
 sg13g2_decap_4 FILLER_40_484 ();
 sg13g2_fill_2 FILLER_40_507 ();
 sg13g2_fill_1 FILLER_40_509 ();
 sg13g2_fill_1 FILLER_40_522 ();
 sg13g2_fill_2 FILLER_40_539 ();
 sg13g2_fill_1 FILLER_40_541 ();
 sg13g2_fill_2 FILLER_40_557 ();
 sg13g2_decap_4 FILLER_40_581 ();
 sg13g2_fill_2 FILLER_40_620 ();
 sg13g2_fill_1 FILLER_40_668 ();
 sg13g2_fill_2 FILLER_40_699 ();
 sg13g2_fill_1 FILLER_40_701 ();
 sg13g2_fill_2 FILLER_40_737 ();
 sg13g2_fill_1 FILLER_40_817 ();
 sg13g2_fill_2 FILLER_40_822 ();
 sg13g2_decap_4 FILLER_40_834 ();
 sg13g2_fill_1 FILLER_40_849 ();
 sg13g2_fill_2 FILLER_40_882 ();
 sg13g2_fill_1 FILLER_40_884 ();
 sg13g2_fill_1 FILLER_40_976 ();
 sg13g2_fill_1 FILLER_40_989 ();
 sg13g2_fill_2 FILLER_40_995 ();
 sg13g2_decap_8 FILLER_41_34 ();
 sg13g2_fill_1 FILLER_41_41 ();
 sg13g2_fill_2 FILLER_41_48 ();
 sg13g2_fill_1 FILLER_41_60 ();
 sg13g2_decap_4 FILLER_41_78 ();
 sg13g2_fill_2 FILLER_41_82 ();
 sg13g2_decap_4 FILLER_41_94 ();
 sg13g2_fill_2 FILLER_41_98 ();
 sg13g2_decap_4 FILLER_41_132 ();
 sg13g2_fill_1 FILLER_41_136 ();
 sg13g2_decap_4 FILLER_41_148 ();
 sg13g2_fill_2 FILLER_41_152 ();
 sg13g2_decap_4 FILLER_41_179 ();
 sg13g2_fill_1 FILLER_41_183 ();
 sg13g2_fill_1 FILLER_41_243 ();
 sg13g2_fill_2 FILLER_41_266 ();
 sg13g2_decap_8 FILLER_41_271 ();
 sg13g2_decap_8 FILLER_41_278 ();
 sg13g2_fill_1 FILLER_41_285 ();
 sg13g2_decap_8 FILLER_41_296 ();
 sg13g2_fill_2 FILLER_41_303 ();
 sg13g2_decap_8 FILLER_41_311 ();
 sg13g2_fill_2 FILLER_41_323 ();
 sg13g2_decap_8 FILLER_41_341 ();
 sg13g2_decap_8 FILLER_41_348 ();
 sg13g2_decap_8 FILLER_41_355 ();
 sg13g2_decap_8 FILLER_41_399 ();
 sg13g2_decap_8 FILLER_41_406 ();
 sg13g2_fill_2 FILLER_41_413 ();
 sg13g2_fill_1 FILLER_41_415 ();
 sg13g2_fill_1 FILLER_41_443 ();
 sg13g2_fill_1 FILLER_41_449 ();
 sg13g2_decap_8 FILLER_41_477 ();
 sg13g2_decap_4 FILLER_41_484 ();
 sg13g2_fill_1 FILLER_41_488 ();
 sg13g2_fill_2 FILLER_41_509 ();
 sg13g2_fill_1 FILLER_41_511 ();
 sg13g2_decap_8 FILLER_41_520 ();
 sg13g2_decap_8 FILLER_41_527 ();
 sg13g2_fill_2 FILLER_41_539 ();
 sg13g2_fill_1 FILLER_41_541 ();
 sg13g2_decap_8 FILLER_41_574 ();
 sg13g2_fill_2 FILLER_41_604 ();
 sg13g2_fill_2 FILLER_41_619 ();
 sg13g2_fill_2 FILLER_41_638 ();
 sg13g2_fill_1 FILLER_41_666 ();
 sg13g2_decap_8 FILLER_41_693 ();
 sg13g2_decap_8 FILLER_41_700 ();
 sg13g2_decap_4 FILLER_41_711 ();
 sg13g2_fill_2 FILLER_41_724 ();
 sg13g2_fill_2 FILLER_41_759 ();
 sg13g2_fill_1 FILLER_41_761 ();
 sg13g2_fill_2 FILLER_41_776 ();
 sg13g2_fill_1 FILLER_41_778 ();
 sg13g2_fill_2 FILLER_41_788 ();
 sg13g2_fill_1 FILLER_41_795 ();
 sg13g2_decap_8 FILLER_41_814 ();
 sg13g2_fill_1 FILLER_41_821 ();
 sg13g2_fill_1 FILLER_41_866 ();
 sg13g2_fill_2 FILLER_41_876 ();
 sg13g2_fill_1 FILLER_41_878 ();
 sg13g2_fill_1 FILLER_41_888 ();
 sg13g2_fill_2 FILLER_41_895 ();
 sg13g2_fill_1 FILLER_41_921 ();
 sg13g2_decap_8 FILLER_41_926 ();
 sg13g2_fill_2 FILLER_41_933 ();
 sg13g2_fill_1 FILLER_41_935 ();
 sg13g2_fill_2 FILLER_41_980 ();
 sg13g2_fill_1 FILLER_41_982 ();
 sg13g2_fill_2 FILLER_41_1001 ();
 sg13g2_decap_4 FILLER_41_1025 ();
 sg13g2_fill_2 FILLER_42_8 ();
 sg13g2_fill_1 FILLER_42_46 ();
 sg13g2_fill_2 FILLER_42_51 ();
 sg13g2_fill_1 FILLER_42_53 ();
 sg13g2_fill_2 FILLER_42_59 ();
 sg13g2_decap_4 FILLER_42_78 ();
 sg13g2_fill_1 FILLER_42_82 ();
 sg13g2_decap_4 FILLER_42_102 ();
 sg13g2_fill_1 FILLER_42_106 ();
 sg13g2_fill_2 FILLER_42_118 ();
 sg13g2_fill_1 FILLER_42_120 ();
 sg13g2_fill_2 FILLER_42_126 ();
 sg13g2_decap_8 FILLER_42_155 ();
 sg13g2_decap_8 FILLER_42_189 ();
 sg13g2_decap_8 FILLER_42_196 ();
 sg13g2_decap_8 FILLER_42_203 ();
 sg13g2_decap_8 FILLER_42_210 ();
 sg13g2_decap_8 FILLER_42_217 ();
 sg13g2_fill_1 FILLER_42_224 ();
 sg13g2_fill_2 FILLER_42_238 ();
 sg13g2_decap_8 FILLER_42_250 ();
 sg13g2_decap_8 FILLER_42_257 ();
 sg13g2_decap_8 FILLER_42_264 ();
 sg13g2_fill_2 FILLER_42_271 ();
 sg13g2_fill_1 FILLER_42_273 ();
 sg13g2_decap_8 FILLER_42_282 ();
 sg13g2_decap_8 FILLER_42_289 ();
 sg13g2_decap_8 FILLER_42_296 ();
 sg13g2_fill_1 FILLER_42_303 ();
 sg13g2_decap_8 FILLER_42_311 ();
 sg13g2_decap_8 FILLER_42_318 ();
 sg13g2_decap_4 FILLER_42_325 ();
 sg13g2_fill_1 FILLER_42_329 ();
 sg13g2_decap_8 FILLER_42_336 ();
 sg13g2_decap_8 FILLER_42_343 ();
 sg13g2_decap_4 FILLER_42_350 ();
 sg13g2_fill_1 FILLER_42_354 ();
 sg13g2_decap_4 FILLER_42_363 ();
 sg13g2_fill_1 FILLER_42_367 ();
 sg13g2_decap_8 FILLER_42_375 ();
 sg13g2_fill_1 FILLER_42_382 ();
 sg13g2_decap_4 FILLER_42_410 ();
 sg13g2_fill_1 FILLER_42_414 ();
 sg13g2_fill_1 FILLER_42_493 ();
 sg13g2_fill_2 FILLER_42_577 ();
 sg13g2_fill_1 FILLER_42_588 ();
 sg13g2_fill_2 FILLER_42_629 ();
 sg13g2_fill_1 FILLER_42_631 ();
 sg13g2_decap_4 FILLER_42_654 ();
 sg13g2_fill_1 FILLER_42_667 ();
 sg13g2_fill_1 FILLER_42_695 ();
 sg13g2_fill_2 FILLER_42_723 ();
 sg13g2_fill_1 FILLER_42_749 ();
 sg13g2_decap_8 FILLER_42_785 ();
 sg13g2_fill_1 FILLER_42_824 ();
 sg13g2_fill_2 FILLER_42_839 ();
 sg13g2_fill_2 FILLER_42_855 ();
 sg13g2_fill_1 FILLER_42_857 ();
 sg13g2_fill_2 FILLER_42_903 ();
 sg13g2_fill_2 FILLER_42_928 ();
 sg13g2_fill_2 FILLER_42_939 ();
 sg13g2_fill_2 FILLER_42_945 ();
 sg13g2_fill_1 FILLER_42_947 ();
 sg13g2_fill_1 FILLER_42_952 ();
 sg13g2_fill_2 FILLER_42_957 ();
 sg13g2_fill_1 FILLER_42_959 ();
 sg13g2_fill_2 FILLER_42_975 ();
 sg13g2_fill_2 FILLER_42_986 ();
 sg13g2_decap_8 FILLER_43_4 ();
 sg13g2_decap_8 FILLER_43_11 ();
 sg13g2_decap_8 FILLER_43_18 ();
 sg13g2_decap_8 FILLER_43_25 ();
 sg13g2_decap_8 FILLER_43_32 ();
 sg13g2_decap_8 FILLER_43_39 ();
 sg13g2_fill_2 FILLER_43_46 ();
 sg13g2_fill_2 FILLER_43_58 ();
 sg13g2_fill_2 FILLER_43_76 ();
 sg13g2_fill_1 FILLER_43_78 ();
 sg13g2_fill_2 FILLER_43_99 ();
 sg13g2_fill_1 FILLER_43_101 ();
 sg13g2_fill_2 FILLER_43_124 ();
 sg13g2_decap_4 FILLER_43_134 ();
 sg13g2_fill_1 FILLER_43_138 ();
 sg13g2_decap_8 FILLER_43_144 ();
 sg13g2_decap_8 FILLER_43_155 ();
 sg13g2_decap_8 FILLER_43_162 ();
 sg13g2_decap_4 FILLER_43_169 ();
 sg13g2_fill_1 FILLER_43_173 ();
 sg13g2_decap_8 FILLER_43_178 ();
 sg13g2_decap_4 FILLER_43_185 ();
 sg13g2_fill_2 FILLER_43_195 ();
 sg13g2_decap_4 FILLER_43_205 ();
 sg13g2_fill_1 FILLER_43_209 ();
 sg13g2_decap_4 FILLER_43_215 ();
 sg13g2_fill_1 FILLER_43_219 ();
 sg13g2_fill_2 FILLER_43_229 ();
 sg13g2_decap_4 FILLER_43_262 ();
 sg13g2_decap_8 FILLER_43_286 ();
 sg13g2_fill_2 FILLER_43_293 ();
 sg13g2_fill_1 FILLER_43_295 ();
 sg13g2_fill_1 FILLER_43_302 ();
 sg13g2_decap_8 FILLER_43_308 ();
 sg13g2_decap_8 FILLER_43_315 ();
 sg13g2_fill_2 FILLER_43_322 ();
 sg13g2_fill_1 FILLER_43_324 ();
 sg13g2_fill_2 FILLER_43_333 ();
 sg13g2_fill_1 FILLER_43_335 ();
 sg13g2_decap_4 FILLER_43_342 ();
 sg13g2_fill_2 FILLER_43_346 ();
 sg13g2_fill_1 FILLER_43_361 ();
 sg13g2_fill_2 FILLER_43_367 ();
 sg13g2_fill_2 FILLER_43_421 ();
 sg13g2_fill_2 FILLER_43_469 ();
 sg13g2_decap_4 FILLER_43_475 ();
 sg13g2_decap_8 FILLER_43_509 ();
 sg13g2_decap_8 FILLER_43_516 ();
 sg13g2_decap_4 FILLER_43_523 ();
 sg13g2_fill_2 FILLER_43_533 ();
 sg13g2_fill_2 FILLER_43_543 ();
 sg13g2_decap_4 FILLER_43_549 ();
 sg13g2_fill_2 FILLER_43_553 ();
 sg13g2_decap_8 FILLER_43_559 ();
 sg13g2_decap_8 FILLER_43_566 ();
 sg13g2_fill_2 FILLER_43_573 ();
 sg13g2_decap_4 FILLER_43_622 ();
 sg13g2_fill_1 FILLER_43_626 ();
 sg13g2_decap_8 FILLER_43_654 ();
 sg13g2_decap_8 FILLER_43_661 ();
 sg13g2_fill_2 FILLER_43_698 ();
 sg13g2_fill_1 FILLER_43_700 ();
 sg13g2_decap_8 FILLER_43_705 ();
 sg13g2_decap_4 FILLER_43_712 ();
 sg13g2_fill_1 FILLER_43_716 ();
 sg13g2_fill_1 FILLER_43_722 ();
 sg13g2_fill_2 FILLER_43_728 ();
 sg13g2_fill_1 FILLER_43_730 ();
 sg13g2_decap_4 FILLER_43_737 ();
 sg13g2_fill_2 FILLER_43_741 ();
 sg13g2_fill_2 FILLER_43_809 ();
 sg13g2_fill_1 FILLER_43_865 ();
 sg13g2_fill_2 FILLER_43_943 ();
 sg13g2_fill_2 FILLER_43_977 ();
 sg13g2_fill_2 FILLER_43_1014 ();
 sg13g2_decap_4 FILLER_43_1025 ();
 sg13g2_fill_2 FILLER_44_4 ();
 sg13g2_fill_1 FILLER_44_6 ();
 sg13g2_decap_8 FILLER_44_32 ();
 sg13g2_fill_2 FILLER_44_39 ();
 sg13g2_fill_2 FILLER_44_88 ();
 sg13g2_fill_2 FILLER_44_108 ();
 sg13g2_fill_2 FILLER_44_120 ();
 sg13g2_decap_4 FILLER_44_138 ();
 sg13g2_decap_4 FILLER_44_148 ();
 sg13g2_fill_2 FILLER_44_152 ();
 sg13g2_decap_4 FILLER_44_159 ();
 sg13g2_fill_1 FILLER_44_163 ();
 sg13g2_decap_4 FILLER_44_194 ();
 sg13g2_decap_8 FILLER_44_253 ();
 sg13g2_fill_1 FILLER_44_260 ();
 sg13g2_decap_4 FILLER_44_281 ();
 sg13g2_fill_2 FILLER_44_312 ();
 sg13g2_fill_1 FILLER_44_314 ();
 sg13g2_decap_4 FILLER_44_335 ();
 sg13g2_decap_8 FILLER_44_370 ();
 sg13g2_decap_4 FILLER_44_377 ();
 sg13g2_fill_1 FILLER_44_381 ();
 sg13g2_decap_4 FILLER_44_471 ();
 sg13g2_fill_2 FILLER_44_475 ();
 sg13g2_fill_1 FILLER_44_494 ();
 sg13g2_decap_8 FILLER_44_511 ();
 sg13g2_decap_4 FILLER_44_518 ();
 sg13g2_fill_1 FILLER_44_522 ();
 sg13g2_decap_4 FILLER_44_552 ();
 sg13g2_fill_2 FILLER_44_562 ();
 sg13g2_fill_1 FILLER_44_564 ();
 sg13g2_decap_8 FILLER_44_569 ();
 sg13g2_fill_2 FILLER_44_576 ();
 sg13g2_fill_2 FILLER_44_583 ();
 sg13g2_fill_1 FILLER_44_606 ();
 sg13g2_decap_4 FILLER_44_652 ();
 sg13g2_fill_1 FILLER_44_656 ();
 sg13g2_decap_4 FILLER_44_709 ();
 sg13g2_fill_2 FILLER_44_740 ();
 sg13g2_fill_1 FILLER_44_742 ();
 sg13g2_fill_1 FILLER_44_762 ();
 sg13g2_fill_1 FILLER_44_772 ();
 sg13g2_decap_4 FILLER_44_782 ();
 sg13g2_fill_2 FILLER_44_786 ();
 sg13g2_fill_1 FILLER_44_850 ();
 sg13g2_decap_4 FILLER_44_927 ();
 sg13g2_fill_1 FILLER_44_931 ();
 sg13g2_decap_8 FILLER_44_937 ();
 sg13g2_decap_4 FILLER_44_944 ();
 sg13g2_fill_2 FILLER_44_948 ();
 sg13g2_decap_4 FILLER_44_954 ();
 sg13g2_fill_1 FILLER_44_958 ();
 sg13g2_fill_1 FILLER_44_969 ();
 sg13g2_fill_2 FILLER_44_988 ();
 sg13g2_fill_2 FILLER_44_1000 ();
 sg13g2_decap_4 FILLER_45_40 ();
 sg13g2_fill_1 FILLER_45_44 ();
 sg13g2_fill_2 FILLER_45_55 ();
 sg13g2_fill_1 FILLER_45_57 ();
 sg13g2_decap_8 FILLER_45_66 ();
 sg13g2_decap_8 FILLER_45_73 ();
 sg13g2_fill_2 FILLER_45_88 ();
 sg13g2_fill_1 FILLER_45_144 ();
 sg13g2_decap_8 FILLER_45_177 ();
 sg13g2_fill_2 FILLER_45_184 ();
 sg13g2_decap_8 FILLER_45_190 ();
 sg13g2_decap_4 FILLER_45_197 ();
 sg13g2_decap_8 FILLER_45_207 ();
 sg13g2_fill_2 FILLER_45_214 ();
 sg13g2_fill_1 FILLER_45_216 ();
 sg13g2_decap_8 FILLER_45_220 ();
 sg13g2_decap_8 FILLER_45_250 ();
 sg13g2_fill_1 FILLER_45_257 ();
 sg13g2_decap_8 FILLER_45_264 ();
 sg13g2_fill_1 FILLER_45_271 ();
 sg13g2_decap_8 FILLER_45_284 ();
 sg13g2_fill_1 FILLER_45_291 ();
 sg13g2_fill_2 FILLER_45_298 ();
 sg13g2_decap_8 FILLER_45_305 ();
 sg13g2_decap_8 FILLER_45_312 ();
 sg13g2_decap_4 FILLER_45_319 ();
 sg13g2_fill_2 FILLER_45_323 ();
 sg13g2_decap_8 FILLER_45_331 ();
 sg13g2_decap_8 FILLER_45_338 ();
 sg13g2_fill_2 FILLER_45_345 ();
 sg13g2_fill_1 FILLER_45_347 ();
 sg13g2_fill_1 FILLER_45_354 ();
 sg13g2_fill_2 FILLER_45_366 ();
 sg13g2_fill_1 FILLER_45_368 ();
 sg13g2_decap_4 FILLER_45_381 ();
 sg13g2_fill_2 FILLER_45_423 ();
 sg13g2_decap_8 FILLER_45_506 ();
 sg13g2_decap_4 FILLER_45_513 ();
 sg13g2_fill_2 FILLER_45_517 ();
 sg13g2_fill_2 FILLER_45_524 ();
 sg13g2_fill_1 FILLER_45_526 ();
 sg13g2_decap_4 FILLER_45_533 ();
 sg13g2_fill_1 FILLER_45_537 ();
 sg13g2_decap_8 FILLER_45_544 ();
 sg13g2_fill_1 FILLER_45_551 ();
 sg13g2_decap_4 FILLER_45_573 ();
 sg13g2_fill_1 FILLER_45_577 ();
 sg13g2_decap_8 FILLER_45_583 ();
 sg13g2_decap_4 FILLER_45_590 ();
 sg13g2_fill_1 FILLER_45_594 ();
 sg13g2_decap_8 FILLER_45_656 ();
 sg13g2_fill_2 FILLER_45_663 ();
 sg13g2_fill_2 FILLER_45_674 ();
 sg13g2_fill_1 FILLER_45_676 ();
 sg13g2_decap_4 FILLER_45_743 ();
 sg13g2_fill_1 FILLER_45_757 ();
 sg13g2_decap_8 FILLER_45_776 ();
 sg13g2_fill_2 FILLER_45_792 ();
 sg13g2_fill_1 FILLER_45_794 ();
 sg13g2_fill_2 FILLER_45_846 ();
 sg13g2_decap_4 FILLER_45_857 ();
 sg13g2_fill_1 FILLER_45_879 ();
 sg13g2_decap_8 FILLER_45_952 ();
 sg13g2_decap_8 FILLER_45_959 ();
 sg13g2_decap_4 FILLER_45_974 ();
 sg13g2_decap_4 FILLER_45_991 ();
 sg13g2_fill_2 FILLER_45_995 ();
 sg13g2_decap_4 FILLER_45_1002 ();
 sg13g2_fill_1 FILLER_45_1006 ();
 sg13g2_decap_8 FILLER_45_1020 ();
 sg13g2_fill_2 FILLER_45_1027 ();
 sg13g2_decap_4 FILLER_46_8 ();
 sg13g2_fill_1 FILLER_46_12 ();
 sg13g2_decap_4 FILLER_46_34 ();
 sg13g2_fill_1 FILLER_46_38 ();
 sg13g2_fill_1 FILLER_46_49 ();
 sg13g2_fill_2 FILLER_46_53 ();
 sg13g2_fill_2 FILLER_46_60 ();
 sg13g2_decap_8 FILLER_46_72 ();
 sg13g2_fill_2 FILLER_46_79 ();
 sg13g2_fill_1 FILLER_46_81 ();
 sg13g2_fill_2 FILLER_46_117 ();
 sg13g2_fill_2 FILLER_46_137 ();
 sg13g2_decap_4 FILLER_46_171 ();
 sg13g2_fill_2 FILLER_46_185 ();
 sg13g2_fill_1 FILLER_46_187 ();
 sg13g2_fill_1 FILLER_46_198 ();
 sg13g2_decap_4 FILLER_46_242 ();
 sg13g2_decap_8 FILLER_46_278 ();
 sg13g2_decap_8 FILLER_46_308 ();
 sg13g2_decap_8 FILLER_46_315 ();
 sg13g2_decap_4 FILLER_46_322 ();
 sg13g2_fill_1 FILLER_46_326 ();
 sg13g2_decap_4 FILLER_46_338 ();
 sg13g2_fill_1 FILLER_46_350 ();
 sg13g2_fill_2 FILLER_46_356 ();
 sg13g2_fill_1 FILLER_46_358 ();
 sg13g2_fill_1 FILLER_46_367 ();
 sg13g2_decap_8 FILLER_46_377 ();
 sg13g2_fill_2 FILLER_46_384 ();
 sg13g2_fill_1 FILLER_46_430 ();
 sg13g2_fill_1 FILLER_46_474 ();
 sg13g2_fill_1 FILLER_46_517 ();
 sg13g2_fill_1 FILLER_46_533 ();
 sg13g2_decap_4 FILLER_46_550 ();
 sg13g2_fill_2 FILLER_46_626 ();
 sg13g2_decap_8 FILLER_46_647 ();
 sg13g2_decap_8 FILLER_46_654 ();
 sg13g2_fill_2 FILLER_46_661 ();
 sg13g2_fill_1 FILLER_46_663 ();
 sg13g2_decap_4 FILLER_46_678 ();
 sg13g2_fill_1 FILLER_46_682 ();
 sg13g2_fill_2 FILLER_46_692 ();
 sg13g2_fill_1 FILLER_46_710 ();
 sg13g2_fill_2 FILLER_46_753 ();
 sg13g2_fill_1 FILLER_46_755 ();
 sg13g2_fill_2 FILLER_46_783 ();
 sg13g2_fill_1 FILLER_46_785 ();
 sg13g2_fill_2 FILLER_46_791 ();
 sg13g2_fill_2 FILLER_46_838 ();
 sg13g2_decap_4 FILLER_46_865 ();
 sg13g2_fill_1 FILLER_46_896 ();
 sg13g2_fill_1 FILLER_46_929 ();
 sg13g2_decap_8 FILLER_46_1021 ();
 sg13g2_fill_1 FILLER_46_1028 ();
 sg13g2_fill_2 FILLER_47_0 ();
 sg13g2_fill_1 FILLER_47_2 ();
 sg13g2_fill_2 FILLER_47_78 ();
 sg13g2_fill_1 FILLER_47_83 ();
 sg13g2_fill_2 FILLER_47_122 ();
 sg13g2_fill_1 FILLER_47_160 ();
 sg13g2_decap_4 FILLER_47_165 ();
 sg13g2_fill_1 FILLER_47_169 ();
 sg13g2_fill_1 FILLER_47_180 ();
 sg13g2_decap_8 FILLER_47_208 ();
 sg13g2_fill_2 FILLER_47_215 ();
 sg13g2_fill_1 FILLER_47_217 ();
 sg13g2_fill_2 FILLER_47_222 ();
 sg13g2_fill_2 FILLER_47_251 ();
 sg13g2_decap_4 FILLER_47_285 ();
 sg13g2_fill_1 FILLER_47_289 ();
 sg13g2_decap_8 FILLER_47_317 ();
 sg13g2_decap_4 FILLER_47_342 ();
 sg13g2_fill_2 FILLER_47_346 ();
 sg13g2_fill_2 FILLER_47_388 ();
 sg13g2_fill_1 FILLER_47_390 ();
 sg13g2_fill_2 FILLER_47_409 ();
 sg13g2_fill_1 FILLER_47_411 ();
 sg13g2_fill_1 FILLER_47_430 ();
 sg13g2_decap_4 FILLER_47_480 ();
 sg13g2_fill_2 FILLER_47_498 ();
 sg13g2_fill_1 FILLER_47_500 ();
 sg13g2_decap_4 FILLER_47_529 ();
 sg13g2_fill_2 FILLER_47_552 ();
 sg13g2_fill_2 FILLER_47_581 ();
 sg13g2_fill_1 FILLER_47_588 ();
 sg13g2_fill_2 FILLER_47_621 ();
 sg13g2_fill_2 FILLER_47_637 ();
 sg13g2_fill_2 FILLER_47_702 ();
 sg13g2_fill_1 FILLER_47_713 ();
 sg13g2_fill_1 FILLER_47_719 ();
 sg13g2_fill_2 FILLER_47_735 ();
 sg13g2_fill_1 FILLER_47_751 ();
 sg13g2_fill_1 FILLER_47_766 ();
 sg13g2_decap_4 FILLER_47_776 ();
 sg13g2_fill_2 FILLER_47_780 ();
 sg13g2_fill_1 FILLER_47_823 ();
 sg13g2_fill_2 FILLER_47_838 ();
 sg13g2_fill_1 FILLER_47_840 ();
 sg13g2_fill_1 FILLER_47_863 ();
 sg13g2_fill_1 FILLER_47_897 ();
 sg13g2_fill_1 FILLER_47_903 ();
 sg13g2_fill_2 FILLER_47_932 ();
 sg13g2_fill_1 FILLER_47_934 ();
 sg13g2_decap_4 FILLER_47_955 ();
 sg13g2_fill_1 FILLER_47_959 ();
 sg13g2_fill_2 FILLER_47_964 ();
 sg13g2_fill_1 FILLER_47_971 ();
 sg13g2_decap_4 FILLER_47_976 ();
 sg13g2_fill_2 FILLER_47_980 ();
 sg13g2_fill_2 FILLER_47_987 ();
 sg13g2_fill_1 FILLER_47_989 ();
 sg13g2_fill_1 FILLER_47_998 ();
 sg13g2_decap_8 FILLER_47_1016 ();
 sg13g2_decap_4 FILLER_47_1023 ();
 sg13g2_fill_2 FILLER_47_1027 ();
 sg13g2_decap_4 FILLER_48_0 ();
 sg13g2_decap_4 FILLER_48_31 ();
 sg13g2_fill_2 FILLER_48_35 ();
 sg13g2_fill_2 FILLER_48_64 ();
 sg13g2_decap_4 FILLER_48_153 ();
 sg13g2_fill_1 FILLER_48_157 ();
 sg13g2_fill_1 FILLER_48_163 ();
 sg13g2_decap_4 FILLER_48_227 ();
 sg13g2_fill_1 FILLER_48_231 ();
 sg13g2_fill_1 FILLER_48_263 ();
 sg13g2_fill_2 FILLER_48_291 ();
 sg13g2_fill_2 FILLER_48_299 ();
 sg13g2_fill_1 FILLER_48_301 ();
 sg13g2_decap_8 FILLER_48_361 ();
 sg13g2_fill_2 FILLER_48_373 ();
 sg13g2_fill_1 FILLER_48_375 ();
 sg13g2_decap_4 FILLER_48_380 ();
 sg13g2_fill_1 FILLER_48_390 ();
 sg13g2_decap_4 FILLER_48_567 ();
 sg13g2_fill_1 FILLER_48_571 ();
 sg13g2_fill_2 FILLER_48_653 ();
 sg13g2_fill_1 FILLER_48_678 ();
 sg13g2_fill_2 FILLER_48_733 ();
 sg13g2_fill_2 FILLER_48_797 ();
 sg13g2_fill_2 FILLER_48_853 ();
 sg13g2_fill_1 FILLER_48_855 ();
 sg13g2_fill_1 FILLER_48_918 ();
 sg13g2_fill_2 FILLER_48_946 ();
 sg13g2_decap_8 FILLER_48_1007 ();
 sg13g2_decap_8 FILLER_48_1014 ();
 sg13g2_decap_8 FILLER_48_1021 ();
 sg13g2_fill_1 FILLER_48_1028 ();
 sg13g2_decap_8 FILLER_49_4 ();
 sg13g2_decap_8 FILLER_49_11 ();
 sg13g2_decap_8 FILLER_49_18 ();
 sg13g2_decap_8 FILLER_49_25 ();
 sg13g2_decap_8 FILLER_49_32 ();
 sg13g2_decap_8 FILLER_49_39 ();
 sg13g2_decap_8 FILLER_49_46 ();
 sg13g2_decap_8 FILLER_49_53 ();
 sg13g2_decap_8 FILLER_49_60 ();
 sg13g2_decap_4 FILLER_49_67 ();
 sg13g2_decap_8 FILLER_49_75 ();
 sg13g2_decap_8 FILLER_49_82 ();
 sg13g2_fill_2 FILLER_49_89 ();
 sg13g2_fill_1 FILLER_49_91 ();
 sg13g2_decap_8 FILLER_49_95 ();
 sg13g2_decap_8 FILLER_49_102 ();
 sg13g2_decap_8 FILLER_49_109 ();
 sg13g2_decap_8 FILLER_49_116 ();
 sg13g2_decap_8 FILLER_49_123 ();
 sg13g2_decap_8 FILLER_49_130 ();
 sg13g2_fill_1 FILLER_49_137 ();
 sg13g2_decap_8 FILLER_49_142 ();
 sg13g2_fill_2 FILLER_49_149 ();
 sg13g2_fill_1 FILLER_49_151 ();
 sg13g2_decap_8 FILLER_49_183 ();
 sg13g2_fill_2 FILLER_49_190 ();
 sg13g2_decap_8 FILLER_49_217 ();
 sg13g2_decap_8 FILLER_49_224 ();
 sg13g2_decap_8 FILLER_49_231 ();
 sg13g2_fill_2 FILLER_49_238 ();
 sg13g2_fill_1 FILLER_49_240 ();
 sg13g2_decap_8 FILLER_49_245 ();
 sg13g2_decap_8 FILLER_49_252 ();
 sg13g2_decap_8 FILLER_49_268 ();
 sg13g2_decap_8 FILLER_49_275 ();
 sg13g2_decap_8 FILLER_49_282 ();
 sg13g2_decap_8 FILLER_49_289 ();
 sg13g2_decap_8 FILLER_49_296 ();
 sg13g2_fill_1 FILLER_49_303 ();
 sg13g2_decap_4 FILLER_49_308 ();
 sg13g2_fill_1 FILLER_49_312 ();
 sg13g2_decap_8 FILLER_49_317 ();
 sg13g2_decap_8 FILLER_49_324 ();
 sg13g2_decap_8 FILLER_49_331 ();
 sg13g2_fill_1 FILLER_49_338 ();
 sg13g2_decap_8 FILLER_49_347 ();
 sg13g2_decap_8 FILLER_49_354 ();
 sg13g2_decap_8 FILLER_49_361 ();
 sg13g2_decap_8 FILLER_49_368 ();
 sg13g2_decap_8 FILLER_49_375 ();
 sg13g2_decap_4 FILLER_49_382 ();
 sg13g2_fill_2 FILLER_49_386 ();
 sg13g2_fill_2 FILLER_49_471 ();
 sg13g2_fill_1 FILLER_49_473 ();
 sg13g2_decap_4 FILLER_49_483 ();
 sg13g2_fill_1 FILLER_49_487 ();
 sg13g2_fill_2 FILLER_49_492 ();
 sg13g2_decap_8 FILLER_49_498 ();
 sg13g2_decap_8 FILLER_49_505 ();
 sg13g2_fill_2 FILLER_49_512 ();
 sg13g2_decap_8 FILLER_49_518 ();
 sg13g2_decap_8 FILLER_49_525 ();
 sg13g2_fill_2 FILLER_49_532 ();
 sg13g2_fill_1 FILLER_49_534 ();
 sg13g2_decap_8 FILLER_49_548 ();
 sg13g2_decap_8 FILLER_49_555 ();
 sg13g2_decap_8 FILLER_49_562 ();
 sg13g2_fill_2 FILLER_49_569 ();
 sg13g2_fill_2 FILLER_49_584 ();
 sg13g2_fill_2 FILLER_49_590 ();
 sg13g2_fill_1 FILLER_49_592 ();
 sg13g2_fill_1 FILLER_49_624 ();
 sg13g2_fill_1 FILLER_49_644 ();
 sg13g2_decap_4 FILLER_49_666 ();
 sg13g2_fill_2 FILLER_49_670 ();
 sg13g2_fill_2 FILLER_49_677 ();
 sg13g2_fill_1 FILLER_49_679 ();
 sg13g2_decap_8 FILLER_49_689 ();
 sg13g2_decap_8 FILLER_49_696 ();
 sg13g2_decap_8 FILLER_49_716 ();
 sg13g2_decap_4 FILLER_49_723 ();
 sg13g2_fill_2 FILLER_49_727 ();
 sg13g2_decap_4 FILLER_49_734 ();
 sg13g2_fill_2 FILLER_49_738 ();
 sg13g2_decap_8 FILLER_49_744 ();
 sg13g2_fill_1 FILLER_49_772 ();
 sg13g2_decap_8 FILLER_49_786 ();
 sg13g2_fill_1 FILLER_49_793 ();
 sg13g2_decap_4 FILLER_49_798 ();
 sg13g2_fill_2 FILLER_49_802 ();
 sg13g2_fill_2 FILLER_49_808 ();
 sg13g2_fill_2 FILLER_49_814 ();
 sg13g2_fill_1 FILLER_49_816 ();
 sg13g2_fill_1 FILLER_49_829 ();
 sg13g2_decap_8 FILLER_49_843 ();
 sg13g2_fill_2 FILLER_49_854 ();
 sg13g2_decap_8 FILLER_49_865 ();
 sg13g2_fill_2 FILLER_49_872 ();
 sg13g2_fill_1 FILLER_49_874 ();
 sg13g2_fill_2 FILLER_49_901 ();
 sg13g2_fill_1 FILLER_49_908 ();
 sg13g2_fill_2 FILLER_49_942 ();
 sg13g2_fill_2 FILLER_49_967 ();
 sg13g2_fill_1 FILLER_49_969 ();
 sg13g2_decap_4 FILLER_49_979 ();
 sg13g2_fill_2 FILLER_49_983 ();
 sg13g2_decap_8 FILLER_49_989 ();
 sg13g2_decap_8 FILLER_49_996 ();
 sg13g2_decap_8 FILLER_49_1003 ();
 sg13g2_decap_8 FILLER_49_1010 ();
 sg13g2_decap_8 FILLER_49_1017 ();
 sg13g2_decap_4 FILLER_49_1024 ();
 sg13g2_fill_1 FILLER_49_1028 ();
endmodule
